// Benchmark "multiplier_sc" written by ABC on Mon Jul 22 15:14:48 2024

module multiplier_sc ( clock, 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0  );
  input  clock;
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0;
  reg lo00, lo01, lo02, lo03, lo04, lo05, lo06, lo07, lo08, lo09, lo10,
    lo11, lo12, lo13, lo14, lo15, lo16, lo17, lo18, lo19, lo20, lo21, lo22,
    lo23, lo24, lo25, lo26, lo27, lo28, lo29, lo30, lo31, lo32, lo33, lo34,
    lo35, lo36, lo37, lo38, lo39, lo40, lo41, lo42, lo43, lo44, lo45, lo46,
    lo47, lo48, lo49, lo50, lo51, lo52, lo53;
  wire new_n178, new_n179, new_n180, new_n182, new_n183, new_n184, new_n185,
    new_n186, new_n187, new_n188, new_n189, new_n190, new_n191, new_n192,
    new_n193, new_n194, new_n195, new_n196, new_n197, new_n198, new_n199,
    new_n200, new_n201, new_n202, new_n203, new_n204, new_n205, new_n206,
    new_n207, new_n208, new_n209, new_n210, new_n211, new_n212, new_n213,
    new_n214, new_n215, new_n216, new_n217, new_n218, new_n219, new_n220,
    new_n221, new_n222, new_n223, new_n224, new_n225, new_n226, new_n227,
    new_n228, new_n229, new_n230, new_n231, new_n232, new_n233, new_n234,
    new_n235, new_n236, new_n237, new_n238, new_n239, new_n240, new_n241,
    new_n242, new_n243, new_n244, new_n245, new_n246, new_n247, new_n248,
    new_n249, new_n250, new_n251, new_n252, new_n253, new_n254, new_n255,
    new_n256, new_n257, new_n258, new_n259, new_n260, new_n261, new_n262,
    new_n263, new_n264, new_n265, new_n266, new_n267, new_n268, new_n269,
    new_n270, new_n271, new_n272, new_n273, new_n274, new_n275, new_n276,
    new_n277, new_n278, new_n279, new_n280, new_n281, new_n282, new_n283,
    new_n284, new_n285, new_n286, new_n287, new_n288, new_n289, new_n290,
    new_n291, new_n292, new_n293, new_n294, new_n295, new_n296, new_n297,
    new_n298, new_n299, new_n300, new_n301, new_n302, new_n303, new_n304,
    new_n305, new_n306, new_n308, new_n309, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n364, new_n365,
    new_n366, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n380, new_n381,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n411, new_n412, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n466, new_n467, new_n468, new_n469,
    new_n470, new_n472, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n479, new_n480, new_n481, new_n482, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n910, new_n912, li00, li01, li02, li03, li04, li05, li06, li07,
    li08, li09, li10, li11, li12, li13, li14, li15, li16, li17, li18, li19,
    li20, li21, li22, li23, li24, li25, li26, li27, li28, li29, li30, li31,
    li32, li33, li34, li35, li36, li37, li38, li39, li40, li41, li42, li43,
    li44, li45, li46, li47, li48, li49, li50, li51, li52, li53;
  assign new_n178 = lo00 & ~lo13;
  assign new_n179 = lo01 & lo13;
  assign new_n180 = ~new_n178 & ~new_n179;
  assign li14 = lo00 & new_n180;
  assign new_n182 = lo00 & ~lo01;
  assign new_n183 = ~lo00 & lo01;
  assign new_n184 = ~new_n182 & ~new_n183;
  assign new_n185 = lo13 & new_n184;
  assign new_n186 = ~lo13 & ~new_n184;
  assign new_n187 = ~new_n185 & ~new_n186;
  assign new_n188 = lo20 & ~lo29;
  assign new_n189 = ~lo20 & lo29;
  assign new_n190 = ~new_n188 & ~new_n189;
  assign new_n191 = lo12 & new_n190;
  assign new_n192 = ~lo12 & ~new_n190;
  assign new_n193 = ~new_n191 & ~new_n192;
  assign new_n194 = lo04 & ~lo07;
  assign new_n195 = ~lo04 & lo07;
  assign new_n196 = ~new_n194 & ~new_n195;
  assign new_n197 = lo03 & ~lo06;
  assign new_n198 = ~lo03 & lo06;
  assign new_n199 = ~new_n197 & ~new_n198;
  assign new_n200 = lo02 & ~lo05;
  assign new_n201 = ~lo02 & lo05;
  assign new_n202 = ~new_n200 & ~new_n201;
  assign new_n203 = new_n199 & new_n202;
  assign new_n204 = new_n196 & new_n203;
  assign new_n205 = lo11 & new_n204;
  assign new_n206 = ~lo11 & ~new_n204;
  assign new_n207 = ~new_n205 & ~new_n206;
  assign new_n208 = ~lo10 & lo53;
  assign new_n209 = lo10 & lo28;
  assign new_n210 = ~new_n208 & ~new_n209;
  assign new_n211 = lo53 & new_n210;
  assign new_n212 = ~lo53 & ~new_n210;
  assign new_n213 = ~new_n211 & ~new_n212;
  assign new_n214 = ~lo10 & lo52;
  assign new_n215 = lo10 & lo27;
  assign new_n216 = ~new_n214 & ~new_n215;
  assign new_n217 = lo52 & new_n216;
  assign new_n218 = ~lo52 & ~new_n216;
  assign new_n219 = ~new_n217 & ~new_n218;
  assign new_n220 = new_n213 & new_n219;
  assign new_n221 = ~lo10 & lo51;
  assign new_n222 = lo10 & lo26;
  assign new_n223 = ~new_n221 & ~new_n222;
  assign new_n224 = lo51 & new_n223;
  assign new_n225 = ~lo51 & ~new_n223;
  assign new_n226 = ~new_n224 & ~new_n225;
  assign new_n227 = ~lo10 & lo50;
  assign new_n228 = lo10 & lo25;
  assign new_n229 = ~new_n227 & ~new_n228;
  assign new_n230 = lo50 & new_n229;
  assign new_n231 = ~lo50 & ~new_n229;
  assign new_n232 = ~new_n230 & ~new_n231;
  assign new_n233 = new_n226 & new_n232;
  assign new_n234 = new_n220 & new_n233;
  assign new_n235 = ~lo10 & lo49;
  assign new_n236 = lo10 & lo24;
  assign new_n237 = ~new_n235 & ~new_n236;
  assign new_n238 = lo49 & new_n237;
  assign new_n239 = ~lo49 & ~new_n237;
  assign new_n240 = ~new_n238 & ~new_n239;
  assign new_n241 = ~lo10 & lo48;
  assign new_n242 = lo10 & lo23;
  assign new_n243 = ~new_n241 & ~new_n242;
  assign new_n244 = lo48 & new_n243;
  assign new_n245 = ~lo48 & ~new_n243;
  assign new_n246 = ~new_n244 & ~new_n245;
  assign new_n247 = new_n240 & new_n246;
  assign new_n248 = ~lo10 & lo47;
  assign new_n249 = lo10 & lo22;
  assign new_n250 = ~new_n248 & ~new_n249;
  assign new_n251 = lo47 & new_n250;
  assign new_n252 = ~lo47 & ~new_n250;
  assign new_n253 = ~new_n251 & ~new_n252;
  assign new_n254 = ~lo10 & lo46;
  assign new_n255 = lo10 & lo21;
  assign new_n256 = ~new_n254 & ~new_n255;
  assign new_n257 = lo46 & new_n256;
  assign new_n258 = ~lo46 & ~new_n256;
  assign new_n259 = ~new_n257 & ~new_n258;
  assign new_n260 = new_n253 & new_n259;
  assign new_n261 = new_n247 & new_n260;
  assign new_n262 = new_n234 & new_n261;
  assign new_n263 = lo10 & new_n262;
  assign new_n264 = ~lo10 & ~new_n262;
  assign new_n265 = ~new_n263 & ~new_n264;
  assign new_n266 = lo33 & ~lo37;
  assign new_n267 = ~lo33 & lo37;
  assign new_n268 = ~new_n266 & ~new_n267;
  assign new_n269 = lo32 & ~lo36;
  assign new_n270 = ~lo32 & lo36;
  assign new_n271 = ~new_n269 & ~new_n270;
  assign new_n272 = new_n268 & new_n271;
  assign new_n273 = lo31 & ~lo35;
  assign new_n274 = ~lo31 & lo35;
  assign new_n275 = ~new_n273 & ~new_n274;
  assign new_n276 = lo30 & ~lo34;
  assign new_n277 = ~lo30 & lo34;
  assign new_n278 = ~new_n276 & ~new_n277;
  assign new_n279 = new_n275 & new_n278;
  assign new_n280 = new_n272 & new_n279;
  assign new_n281 = lo09 & new_n280;
  assign new_n282 = ~lo09 & ~new_n280;
  assign new_n283 = ~new_n281 & ~new_n282;
  assign new_n284 = lo41 & ~lo45;
  assign new_n285 = ~lo41 & lo45;
  assign new_n286 = ~new_n284 & ~new_n285;
  assign new_n287 = lo40 & ~lo44;
  assign new_n288 = ~lo40 & lo44;
  assign new_n289 = ~new_n287 & ~new_n288;
  assign new_n290 = new_n286 & new_n289;
  assign new_n291 = lo39 & ~lo43;
  assign new_n292 = ~lo39 & lo43;
  assign new_n293 = ~new_n291 & ~new_n292;
  assign new_n294 = lo38 & ~lo42;
  assign new_n295 = ~lo38 & lo42;
  assign new_n296 = ~new_n294 & ~new_n295;
  assign new_n297 = new_n293 & new_n296;
  assign new_n298 = new_n290 & new_n297;
  assign new_n299 = lo08 & new_n298;
  assign new_n300 = ~lo08 & ~new_n298;
  assign new_n301 = ~new_n299 & ~new_n300;
  assign new_n302 = ~lo19 & new_n301;
  assign new_n303 = new_n283 & new_n302;
  assign new_n304 = new_n265 & new_n303;
  assign new_n305 = new_n207 & new_n304;
  assign new_n306 = new_n193 & new_n305;
  assign li19 = ~new_n187 | ~new_n306;
  assign new_n308 = lo00 & ~new_n262;
  assign new_n309 = ~new_n180 & new_n308;
  assign li17 = lo17 | new_n309;
  assign new_n311 = ~li19 & ~li17;
  assign new_n312 = ~li14 & new_n311;
  assign new_n313 = lo00 & ~new_n312;
  assign new_n314 = ~lo32 & ~lo33;
  assign new_n315 = ~lo30 & ~lo31;
  assign new_n316 = new_n314 & new_n315;
  assign new_n317 = ~lo40 & ~lo41;
  assign new_n318 = ~lo38 & ~lo39;
  assign new_n319 = new_n317 & new_n318;
  assign new_n320 = ~new_n316 & ~new_n319;
  assign new_n321 = lo20 & ~new_n320;
  assign new_n322 = new_n312 & new_n321;
  assign li00 = new_n313 | new_n322;
  assign li15 = ~lo00 & ~new_n180;
  assign new_n325 = new_n311 & ~li15;
  assign new_n326 = ~new_n180 & ~new_n325;
  assign new_n327 = ~lo09 & lo32;
  assign new_n328 = lo09 & lo36;
  assign new_n329 = ~new_n327 & ~new_n328;
  assign new_n330 = ~lo09 & lo33;
  assign new_n331 = lo09 & lo37;
  assign new_n332 = ~new_n330 & ~new_n331;
  assign new_n333 = new_n329 & new_n332;
  assign new_n334 = ~lo09 & lo31;
  assign new_n335 = lo09 & lo35;
  assign new_n336 = ~new_n334 & ~new_n335;
  assign new_n337 = ~lo09 & lo30;
  assign new_n338 = lo09 & lo34;
  assign new_n339 = ~new_n337 & ~new_n338;
  assign new_n340 = new_n336 & new_n339;
  assign new_n341 = new_n333 & new_n340;
  assign new_n342 = ~lo08 & lo40;
  assign new_n343 = lo08 & lo44;
  assign new_n344 = ~new_n342 & ~new_n343;
  assign new_n345 = ~lo08 & lo41;
  assign new_n346 = lo08 & lo45;
  assign new_n347 = ~new_n345 & ~new_n346;
  assign new_n348 = new_n344 & new_n347;
  assign new_n349 = ~lo08 & lo38;
  assign new_n350 = lo08 & lo42;
  assign new_n351 = ~new_n349 & ~new_n350;
  assign new_n352 = ~lo08 & lo39;
  assign new_n353 = lo08 & lo43;
  assign new_n354 = ~new_n352 & ~new_n353;
  assign new_n355 = new_n351 & new_n354;
  assign new_n356 = new_n348 & new_n355;
  assign new_n357 = ~new_n341 & ~new_n356;
  assign new_n358 = ~lo12 & lo20;
  assign new_n359 = lo12 & lo29;
  assign new_n360 = ~new_n358 & ~new_n359;
  assign new_n361 = ~new_n357 & ~new_n360;
  assign new_n362 = new_n325 & new_n361;
  assign li01 = new_n326 | new_n362;
  assign new_n364 = lo02 & ~new_n312;
  assign new_n365 = ~lo02 & lo20;
  assign new_n366 = new_n312 & new_n365;
  assign li02 = new_n364 | new_n366;
  assign new_n368 = lo03 & ~new_n312;
  assign new_n369 = ~lo02 & lo03;
  assign new_n370 = lo02 & ~lo03;
  assign new_n371 = ~new_n369 & ~new_n370;
  assign new_n372 = lo20 & ~new_n371;
  assign new_n373 = new_n312 & new_n372;
  assign li03 = new_n368 | new_n373;
  assign new_n375 = lo04 & ~new_n312;
  assign new_n376 = lo02 & lo03;
  assign new_n377 = lo04 & ~new_n376;
  assign new_n378 = ~lo04 & new_n376;
  assign new_n379 = ~new_n377 & ~new_n378;
  assign new_n380 = lo20 & ~new_n379;
  assign new_n381 = new_n312 & new_n380;
  assign li04 = new_n375 | new_n381;
  assign new_n383 = lo02 & ~lo11;
  assign new_n384 = lo05 & lo11;
  assign new_n385 = ~new_n383 & ~new_n384;
  assign new_n386 = ~new_n325 & ~new_n385;
  assign new_n387 = ~new_n360 & new_n385;
  assign new_n388 = new_n325 & new_n387;
  assign li05 = new_n386 | new_n388;
  assign new_n390 = lo03 & ~lo11;
  assign new_n391 = lo06 & lo11;
  assign new_n392 = ~new_n390 & ~new_n391;
  assign new_n393 = ~new_n325 & ~new_n392;
  assign new_n394 = new_n385 & ~new_n392;
  assign new_n395 = ~new_n385 & new_n392;
  assign new_n396 = ~new_n394 & ~new_n395;
  assign new_n397 = ~new_n360 & ~new_n396;
  assign new_n398 = new_n325 & new_n397;
  assign li06 = new_n393 | new_n398;
  assign new_n400 = lo04 & ~lo11;
  assign new_n401 = lo07 & lo11;
  assign new_n402 = ~new_n400 & ~new_n401;
  assign new_n403 = ~new_n325 & ~new_n402;
  assign new_n404 = ~new_n385 & ~new_n392;
  assign new_n405 = ~new_n402 & ~new_n404;
  assign new_n406 = new_n402 & new_n404;
  assign new_n407 = ~new_n405 & ~new_n406;
  assign new_n408 = ~new_n360 & ~new_n407;
  assign new_n409 = new_n325 & new_n408;
  assign li07 = new_n403 | new_n409;
  assign new_n411 = lo08 & ~new_n311;
  assign new_n412 = ~new_n325 & ~new_n347;
  assign new_n413 = pi13 & new_n360;
  assign new_n414 = pi08 & new_n413;
  assign new_n415 = ~new_n347 & ~new_n413;
  assign new_n416 = ~new_n414 & ~new_n415;
  assign new_n417 = new_n325 & ~new_n416;
  assign li45 = new_n412 | new_n417;
  assign new_n419 = lo41 & ~new_n312;
  assign new_n420 = pi13 & ~lo20;
  assign new_n421 = pi04 & new_n420;
  assign new_n422 = lo41 & ~new_n420;
  assign new_n423 = ~new_n421 & ~new_n422;
  assign new_n424 = new_n312 & ~new_n423;
  assign li41 = new_n419 | new_n424;
  assign new_n426 = ~li45 & li41;
  assign new_n427 = li45 & ~li41;
  assign new_n428 = ~new_n426 & ~new_n427;
  assign new_n429 = ~new_n325 & ~new_n344;
  assign new_n430 = pi07 & new_n413;
  assign new_n431 = ~new_n344 & ~new_n413;
  assign new_n432 = ~new_n430 & ~new_n431;
  assign new_n433 = new_n325 & ~new_n432;
  assign li44 = new_n429 | new_n433;
  assign new_n435 = lo40 & ~new_n312;
  assign new_n436 = pi03 & new_n420;
  assign new_n437 = lo40 & ~new_n420;
  assign new_n438 = ~new_n436 & ~new_n437;
  assign new_n439 = new_n312 & ~new_n438;
  assign li40 = new_n435 | new_n439;
  assign new_n441 = ~li44 & li40;
  assign new_n442 = li44 & ~li40;
  assign new_n443 = ~new_n441 & ~new_n442;
  assign new_n444 = new_n428 & new_n443;
  assign new_n445 = ~new_n325 & ~new_n354;
  assign new_n446 = pi06 & new_n413;
  assign new_n447 = ~new_n354 & ~new_n413;
  assign new_n448 = ~new_n446 & ~new_n447;
  assign new_n449 = new_n325 & ~new_n448;
  assign li43 = new_n445 | new_n449;
  assign new_n451 = lo39 & ~new_n312;
  assign new_n452 = pi02 & new_n420;
  assign new_n453 = lo39 & ~new_n420;
  assign new_n454 = ~new_n452 & ~new_n453;
  assign new_n455 = new_n312 & ~new_n454;
  assign li39 = new_n451 | new_n455;
  assign new_n457 = ~li43 & li39;
  assign new_n458 = li43 & ~li39;
  assign new_n459 = ~new_n457 & ~new_n458;
  assign new_n460 = ~new_n325 & ~new_n351;
  assign new_n461 = pi05 & new_n413;
  assign new_n462 = ~new_n351 & ~new_n413;
  assign new_n463 = ~new_n461 & ~new_n462;
  assign new_n464 = new_n325 & ~new_n463;
  assign li42 = new_n460 | new_n464;
  assign new_n466 = lo38 & ~new_n312;
  assign new_n467 = pi01 & new_n420;
  assign new_n468 = lo38 & ~new_n420;
  assign new_n469 = ~new_n467 & ~new_n468;
  assign new_n470 = new_n312 & ~new_n469;
  assign li38 = new_n466 | new_n470;
  assign new_n472 = ~li42 & li38;
  assign new_n473 = li42 & ~li38;
  assign new_n474 = ~new_n472 & ~new_n473;
  assign new_n475 = new_n459 & new_n474;
  assign new_n476 = new_n444 & new_n475;
  assign new_n477 = new_n311 & ~new_n476;
  assign li08 = new_n411 | new_n477;
  assign new_n479 = lo09 & ~new_n311;
  assign new_n480 = ~new_n325 & ~new_n332;
  assign new_n481 = pi12 & new_n413;
  assign new_n482 = new_n325 & new_n481;
  assign li37 = new_n480 | new_n482;
  assign new_n484 = lo33 & ~new_n312;
  assign new_n485 = pi12 & new_n420;
  assign new_n486 = new_n312 & new_n485;
  assign li33 = new_n484 | new_n486;
  assign new_n488 = ~li37 & li33;
  assign new_n489 = li37 & ~li33;
  assign new_n490 = ~new_n488 & ~new_n489;
  assign new_n491 = ~new_n325 & ~new_n329;
  assign new_n492 = pi11 & new_n413;
  assign new_n493 = ~new_n332 & ~new_n413;
  assign new_n494 = ~new_n492 & ~new_n493;
  assign new_n495 = new_n325 & ~new_n494;
  assign li36 = new_n491 | new_n495;
  assign new_n497 = lo32 & ~new_n312;
  assign new_n498 = pi11 & new_n420;
  assign new_n499 = lo33 & ~new_n420;
  assign new_n500 = ~new_n498 & ~new_n499;
  assign new_n501 = new_n312 & ~new_n500;
  assign li32 = new_n497 | new_n501;
  assign new_n503 = ~li36 & li32;
  assign new_n504 = li36 & ~li32;
  assign new_n505 = ~new_n503 & ~new_n504;
  assign new_n506 = new_n490 & new_n505;
  assign new_n507 = ~new_n325 & ~new_n336;
  assign new_n508 = pi10 & new_n413;
  assign new_n509 = ~new_n329 & ~new_n413;
  assign new_n510 = ~new_n508 & ~new_n509;
  assign new_n511 = new_n325 & ~new_n510;
  assign li35 = new_n507 | new_n511;
  assign new_n513 = lo31 & ~new_n312;
  assign new_n514 = pi10 & new_n420;
  assign new_n515 = lo32 & ~new_n420;
  assign new_n516 = ~new_n514 & ~new_n515;
  assign new_n517 = new_n312 & ~new_n516;
  assign li31 = new_n513 | new_n517;
  assign new_n519 = ~li35 & li31;
  assign new_n520 = li35 & ~li31;
  assign new_n521 = ~new_n519 & ~new_n520;
  assign new_n522 = ~new_n325 & ~new_n339;
  assign new_n523 = pi09 & new_n413;
  assign new_n524 = ~new_n336 & ~new_n413;
  assign new_n525 = ~new_n523 & ~new_n524;
  assign new_n526 = new_n325 & ~new_n525;
  assign li34 = new_n522 | new_n526;
  assign new_n528 = lo30 & ~new_n312;
  assign new_n529 = pi09 & new_n420;
  assign new_n530 = lo31 & ~new_n420;
  assign new_n531 = ~new_n529 & ~new_n530;
  assign new_n532 = new_n312 & ~new_n531;
  assign li30 = new_n528 | new_n532;
  assign new_n534 = ~li34 & li30;
  assign new_n535 = li34 & ~li30;
  assign new_n536 = ~new_n534 & ~new_n535;
  assign new_n537 = new_n521 & new_n536;
  assign new_n538 = new_n506 & new_n537;
  assign new_n539 = new_n311 & ~new_n538;
  assign li09 = new_n479 | new_n539;
  assign new_n541 = lo10 & ~new_n311;
  assign new_n542 = ~new_n210 & ~new_n325;
  assign new_n543 = ~new_n351 & new_n385;
  assign new_n544 = new_n392 & new_n543;
  assign new_n545 = new_n402 & new_n544;
  assign new_n546 = ~new_n339 & new_n545;
  assign new_n547 = ~new_n256 & new_n546;
  assign new_n548 = ~new_n351 & ~new_n385;
  assign new_n549 = ~new_n354 & new_n385;
  assign new_n550 = ~new_n548 & ~new_n549;
  assign new_n551 = new_n392 & ~new_n550;
  assign new_n552 = new_n402 & new_n551;
  assign new_n553 = ~new_n339 & new_n552;
  assign new_n554 = new_n250 & new_n553;
  assign new_n555 = ~new_n250 & ~new_n553;
  assign new_n556 = ~new_n554 & ~new_n555;
  assign new_n557 = new_n547 & ~new_n556;
  assign new_n558 = ~new_n250 & new_n553;
  assign new_n559 = ~new_n557 & ~new_n558;
  assign new_n560 = ~new_n392 & new_n543;
  assign new_n561 = ~new_n354 & ~new_n385;
  assign new_n562 = ~new_n344 & new_n385;
  assign new_n563 = ~new_n561 & ~new_n562;
  assign new_n564 = new_n392 & ~new_n563;
  assign new_n565 = ~new_n560 & ~new_n564;
  assign new_n566 = new_n402 & ~new_n565;
  assign new_n567 = ~new_n339 & new_n566;
  assign new_n568 = new_n243 & new_n567;
  assign new_n569 = ~new_n243 & ~new_n567;
  assign new_n570 = ~new_n568 & ~new_n569;
  assign new_n571 = ~new_n392 & ~new_n550;
  assign new_n572 = ~new_n344 & ~new_n385;
  assign new_n573 = ~new_n347 & new_n385;
  assign new_n574 = ~new_n572 & ~new_n573;
  assign new_n575 = new_n392 & ~new_n574;
  assign new_n576 = ~new_n571 & ~new_n575;
  assign new_n577 = new_n402 & ~new_n576;
  assign new_n578 = ~new_n339 & new_n577;
  assign new_n579 = new_n237 & new_n578;
  assign new_n580 = ~new_n237 & ~new_n578;
  assign new_n581 = ~new_n579 & ~new_n580;
  assign new_n582 = ~new_n570 & ~new_n581;
  assign new_n583 = ~new_n559 & new_n582;
  assign new_n584 = ~new_n243 & new_n567;
  assign new_n585 = ~new_n581 & new_n584;
  assign new_n586 = ~new_n237 & new_n578;
  assign new_n587 = ~new_n585 & ~new_n586;
  assign new_n588 = ~new_n583 & new_n587;
  assign new_n589 = ~new_n402 & new_n544;
  assign new_n590 = ~new_n392 & ~new_n563;
  assign new_n591 = ~new_n347 & ~new_n385;
  assign new_n592 = new_n392 & new_n591;
  assign new_n593 = ~new_n590 & ~new_n592;
  assign new_n594 = new_n402 & ~new_n593;
  assign new_n595 = ~new_n589 & ~new_n594;
  assign new_n596 = ~new_n339 & ~new_n595;
  assign new_n597 = new_n229 & new_n596;
  assign new_n598 = ~new_n229 & ~new_n596;
  assign new_n599 = ~new_n597 & ~new_n598;
  assign new_n600 = ~new_n402 & new_n551;
  assign new_n601 = ~new_n392 & ~new_n574;
  assign new_n602 = new_n402 & new_n601;
  assign new_n603 = ~new_n600 & ~new_n602;
  assign new_n604 = ~new_n339 & ~new_n603;
  assign new_n605 = new_n223 & new_n604;
  assign new_n606 = ~new_n223 & ~new_n604;
  assign new_n607 = ~new_n605 & ~new_n606;
  assign new_n608 = ~new_n599 & ~new_n607;
  assign new_n609 = ~new_n588 & new_n608;
  assign new_n610 = ~new_n229 & new_n596;
  assign new_n611 = ~new_n607 & new_n610;
  assign new_n612 = ~new_n223 & new_n604;
  assign new_n613 = ~new_n611 & ~new_n612;
  assign new_n614 = ~new_n609 & new_n613;
  assign new_n615 = ~new_n402 & ~new_n565;
  assign new_n616 = ~new_n392 & new_n591;
  assign new_n617 = new_n402 & new_n616;
  assign new_n618 = ~new_n615 & ~new_n617;
  assign new_n619 = ~new_n339 & ~new_n618;
  assign new_n620 = new_n216 & new_n619;
  assign new_n621 = ~new_n216 & ~new_n619;
  assign new_n622 = ~new_n620 & ~new_n621;
  assign new_n623 = ~new_n614 & ~new_n622;
  assign new_n624 = ~new_n216 & new_n619;
  assign new_n625 = ~new_n623 & ~new_n624;
  assign new_n626 = ~new_n402 & ~new_n576;
  assign new_n627 = ~new_n339 & new_n626;
  assign new_n628 = new_n210 & new_n627;
  assign new_n629 = ~new_n210 & ~new_n627;
  assign new_n630 = ~new_n628 & ~new_n629;
  assign new_n631 = new_n625 & ~new_n630;
  assign new_n632 = ~new_n625 & new_n630;
  assign new_n633 = ~new_n631 & ~new_n632;
  assign new_n634 = ~new_n360 & ~new_n633;
  assign new_n635 = new_n325 & new_n634;
  assign li28 = new_n542 | new_n635;
  assign new_n637 = lo53 & ~new_n312;
  assign new_n638 = ~lo02 & lo38;
  assign new_n639 = ~lo03 & new_n638;
  assign new_n640 = ~lo04 & new_n639;
  assign new_n641 = lo30 & new_n640;
  assign new_n642 = lo46 & new_n641;
  assign new_n643 = lo02 & lo38;
  assign new_n644 = ~lo02 & lo39;
  assign new_n645 = ~new_n643 & ~new_n644;
  assign new_n646 = ~lo03 & ~new_n645;
  assign new_n647 = ~lo04 & new_n646;
  assign new_n648 = lo30 & new_n647;
  assign new_n649 = ~lo47 & new_n648;
  assign new_n650 = lo47 & ~new_n648;
  assign new_n651 = ~new_n649 & ~new_n650;
  assign new_n652 = new_n642 & ~new_n651;
  assign new_n653 = lo47 & new_n648;
  assign new_n654 = ~new_n652 & ~new_n653;
  assign new_n655 = lo03 & new_n638;
  assign new_n656 = lo02 & lo39;
  assign new_n657 = ~lo02 & lo40;
  assign new_n658 = ~new_n656 & ~new_n657;
  assign new_n659 = ~lo03 & ~new_n658;
  assign new_n660 = ~new_n655 & ~new_n659;
  assign new_n661 = ~lo04 & ~new_n660;
  assign new_n662 = lo30 & new_n661;
  assign new_n663 = ~lo48 & new_n662;
  assign new_n664 = lo48 & ~new_n662;
  assign new_n665 = ~new_n663 & ~new_n664;
  assign new_n666 = lo03 & ~new_n645;
  assign new_n667 = lo02 & lo40;
  assign new_n668 = ~lo02 & lo41;
  assign new_n669 = ~new_n667 & ~new_n668;
  assign new_n670 = ~lo03 & ~new_n669;
  assign new_n671 = ~new_n666 & ~new_n670;
  assign new_n672 = ~lo04 & ~new_n671;
  assign new_n673 = lo30 & new_n672;
  assign new_n674 = ~lo49 & new_n673;
  assign new_n675 = lo49 & ~new_n673;
  assign new_n676 = ~new_n674 & ~new_n675;
  assign new_n677 = ~new_n665 & ~new_n676;
  assign new_n678 = ~new_n654 & new_n677;
  assign new_n679 = lo48 & new_n662;
  assign new_n680 = ~new_n676 & new_n679;
  assign new_n681 = lo49 & new_n673;
  assign new_n682 = ~new_n680 & ~new_n681;
  assign new_n683 = ~new_n678 & new_n682;
  assign new_n684 = lo04 & new_n639;
  assign new_n685 = lo03 & ~new_n658;
  assign new_n686 = lo02 & lo41;
  assign new_n687 = ~lo03 & new_n686;
  assign new_n688 = ~new_n685 & ~new_n687;
  assign new_n689 = ~lo04 & ~new_n688;
  assign new_n690 = ~new_n684 & ~new_n689;
  assign new_n691 = lo30 & ~new_n690;
  assign new_n692 = ~lo50 & new_n691;
  assign new_n693 = lo50 & ~new_n691;
  assign new_n694 = ~new_n692 & ~new_n693;
  assign new_n695 = lo04 & new_n646;
  assign new_n696 = lo03 & ~new_n669;
  assign new_n697 = ~lo04 & new_n696;
  assign new_n698 = ~new_n695 & ~new_n697;
  assign new_n699 = lo30 & ~new_n698;
  assign new_n700 = ~lo51 & new_n699;
  assign new_n701 = lo51 & ~new_n699;
  assign new_n702 = ~new_n700 & ~new_n701;
  assign new_n703 = ~new_n694 & ~new_n702;
  assign new_n704 = ~new_n683 & new_n703;
  assign new_n705 = lo50 & new_n691;
  assign new_n706 = ~new_n702 & new_n705;
  assign new_n707 = lo51 & new_n699;
  assign new_n708 = ~new_n706 & ~new_n707;
  assign new_n709 = ~new_n704 & new_n708;
  assign new_n710 = lo04 & ~new_n660;
  assign new_n711 = lo03 & new_n686;
  assign new_n712 = ~lo04 & new_n711;
  assign new_n713 = ~new_n710 & ~new_n712;
  assign new_n714 = lo30 & ~new_n713;
  assign new_n715 = ~lo52 & new_n714;
  assign new_n716 = lo52 & ~new_n714;
  assign new_n717 = ~new_n715 & ~new_n716;
  assign new_n718 = ~new_n709 & ~new_n717;
  assign new_n719 = lo52 & new_n714;
  assign new_n720 = ~new_n718 & ~new_n719;
  assign new_n721 = lo04 & ~new_n671;
  assign new_n722 = lo30 & new_n721;
  assign new_n723 = ~lo53 & new_n722;
  assign new_n724 = lo53 & ~new_n722;
  assign new_n725 = ~new_n723 & ~new_n724;
  assign new_n726 = new_n720 & ~new_n725;
  assign new_n727 = ~new_n720 & new_n725;
  assign new_n728 = ~new_n726 & ~new_n727;
  assign new_n729 = lo20 & ~new_n728;
  assign new_n730 = new_n312 & new_n729;
  assign li53 = new_n637 | new_n730;
  assign new_n732 = ~li28 & li53;
  assign new_n733 = li28 & ~li53;
  assign new_n734 = ~new_n732 & ~new_n733;
  assign new_n735 = ~new_n216 & ~new_n325;
  assign new_n736 = new_n614 & ~new_n622;
  assign new_n737 = ~new_n614 & new_n622;
  assign new_n738 = ~new_n736 & ~new_n737;
  assign new_n739 = ~new_n360 & ~new_n738;
  assign new_n740 = new_n325 & new_n739;
  assign li27 = new_n735 | new_n740;
  assign new_n742 = lo52 & ~new_n312;
  assign new_n743 = new_n709 & ~new_n717;
  assign new_n744 = ~new_n709 & new_n717;
  assign new_n745 = ~new_n743 & ~new_n744;
  assign new_n746 = lo20 & ~new_n745;
  assign new_n747 = new_n312 & new_n746;
  assign li52 = new_n742 | new_n747;
  assign new_n749 = ~li27 & li52;
  assign new_n750 = li27 & ~li52;
  assign new_n751 = ~new_n749 & ~new_n750;
  assign new_n752 = new_n734 & new_n751;
  assign new_n753 = ~new_n223 & ~new_n325;
  assign new_n754 = ~new_n588 & ~new_n599;
  assign new_n755 = ~new_n610 & ~new_n754;
  assign new_n756 = ~new_n607 & new_n755;
  assign new_n757 = new_n607 & ~new_n755;
  assign new_n758 = ~new_n756 & ~new_n757;
  assign new_n759 = ~new_n360 & ~new_n758;
  assign new_n760 = new_n325 & new_n759;
  assign li26 = new_n753 | new_n760;
  assign new_n762 = lo51 & ~new_n312;
  assign new_n763 = ~new_n683 & ~new_n694;
  assign new_n764 = ~new_n705 & ~new_n763;
  assign new_n765 = ~new_n702 & new_n764;
  assign new_n766 = new_n702 & ~new_n764;
  assign new_n767 = ~new_n765 & ~new_n766;
  assign new_n768 = lo20 & ~new_n767;
  assign new_n769 = new_n312 & new_n768;
  assign li51 = new_n762 | new_n769;
  assign new_n771 = ~li26 & li51;
  assign new_n772 = li26 & ~li51;
  assign new_n773 = ~new_n771 & ~new_n772;
  assign new_n774 = ~new_n229 & ~new_n325;
  assign new_n775 = new_n588 & ~new_n599;
  assign new_n776 = ~new_n588 & new_n599;
  assign new_n777 = ~new_n775 & ~new_n776;
  assign new_n778 = ~new_n360 & ~new_n777;
  assign new_n779 = new_n325 & new_n778;
  assign li25 = new_n774 | new_n779;
  assign new_n781 = lo50 & ~new_n312;
  assign new_n782 = new_n683 & ~new_n694;
  assign new_n783 = ~new_n683 & new_n694;
  assign new_n784 = ~new_n782 & ~new_n783;
  assign new_n785 = lo20 & ~new_n784;
  assign new_n786 = new_n312 & new_n785;
  assign li50 = new_n781 | new_n786;
  assign new_n788 = ~li25 & li50;
  assign new_n789 = li25 & ~li50;
  assign new_n790 = ~new_n788 & ~new_n789;
  assign new_n791 = new_n773 & new_n790;
  assign new_n792 = new_n752 & new_n791;
  assign new_n793 = ~new_n237 & ~new_n325;
  assign new_n794 = ~new_n559 & ~new_n570;
  assign new_n795 = ~new_n584 & ~new_n794;
  assign new_n796 = ~new_n581 & new_n795;
  assign new_n797 = new_n581 & ~new_n795;
  assign new_n798 = ~new_n796 & ~new_n797;
  assign new_n799 = ~new_n360 & ~new_n798;
  assign new_n800 = new_n325 & new_n799;
  assign li24 = new_n793 | new_n800;
  assign new_n802 = lo49 & ~new_n312;
  assign new_n803 = ~new_n654 & ~new_n665;
  assign new_n804 = ~new_n679 & ~new_n803;
  assign new_n805 = ~new_n676 & new_n804;
  assign new_n806 = new_n676 & ~new_n804;
  assign new_n807 = ~new_n805 & ~new_n806;
  assign new_n808 = lo20 & ~new_n807;
  assign new_n809 = new_n312 & new_n808;
  assign li49 = new_n802 | new_n809;
  assign new_n811 = ~li24 & li49;
  assign new_n812 = li24 & ~li49;
  assign new_n813 = ~new_n811 & ~new_n812;
  assign new_n814 = ~new_n243 & ~new_n325;
  assign new_n815 = new_n559 & ~new_n570;
  assign new_n816 = ~new_n559 & new_n570;
  assign new_n817 = ~new_n815 & ~new_n816;
  assign new_n818 = ~new_n360 & ~new_n817;
  assign new_n819 = new_n325 & new_n818;
  assign li23 = new_n814 | new_n819;
  assign new_n821 = lo48 & ~new_n312;
  assign new_n822 = new_n654 & ~new_n665;
  assign new_n823 = ~new_n654 & new_n665;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = lo20 & ~new_n824;
  assign new_n826 = new_n312 & new_n825;
  assign li48 = new_n821 | new_n826;
  assign new_n828 = ~li23 & li48;
  assign new_n829 = li23 & ~li48;
  assign new_n830 = ~new_n828 & ~new_n829;
  assign new_n831 = new_n813 & new_n830;
  assign new_n832 = ~new_n250 & ~new_n325;
  assign new_n833 = ~new_n547 & ~new_n556;
  assign new_n834 = new_n547 & new_n556;
  assign new_n835 = ~new_n833 & ~new_n834;
  assign new_n836 = ~new_n360 & ~new_n835;
  assign new_n837 = new_n325 & new_n836;
  assign li22 = new_n832 | new_n837;
  assign new_n839 = lo47 & ~new_n312;
  assign new_n840 = ~new_n642 & ~new_n651;
  assign new_n841 = new_n642 & new_n651;
  assign new_n842 = ~new_n840 & ~new_n841;
  assign new_n843 = lo20 & ~new_n842;
  assign new_n844 = new_n312 & new_n843;
  assign li47 = new_n839 | new_n844;
  assign new_n846 = ~li22 & li47;
  assign new_n847 = li22 & ~li47;
  assign new_n848 = ~new_n846 & ~new_n847;
  assign new_n849 = ~new_n256 & ~new_n325;
  assign new_n850 = new_n256 & new_n546;
  assign new_n851 = ~new_n256 & ~new_n546;
  assign new_n852 = ~new_n850 & ~new_n851;
  assign new_n853 = ~new_n360 & ~new_n852;
  assign new_n854 = new_n325 & new_n853;
  assign li21 = new_n849 | new_n854;
  assign new_n856 = lo46 & ~new_n312;
  assign new_n857 = ~lo46 & new_n641;
  assign new_n858 = lo46 & ~new_n641;
  assign new_n859 = ~new_n857 & ~new_n858;
  assign new_n860 = lo20 & ~new_n859;
  assign new_n861 = new_n312 & new_n860;
  assign li46 = new_n856 | new_n861;
  assign new_n863 = ~li21 & li46;
  assign new_n864 = li21 & ~li46;
  assign new_n865 = ~new_n863 & ~new_n864;
  assign new_n866 = new_n848 & new_n865;
  assign new_n867 = new_n831 & new_n866;
  assign new_n868 = new_n792 & new_n867;
  assign new_n869 = new_n311 & ~new_n868;
  assign li10 = new_n541 | new_n869;
  assign new_n871 = lo11 & ~new_n311;
  assign new_n872 = li04 & ~li07;
  assign new_n873 = ~li04 & li07;
  assign new_n874 = ~new_n872 & ~new_n873;
  assign new_n875 = li03 & ~li06;
  assign new_n876 = ~li03 & li06;
  assign new_n877 = ~new_n875 & ~new_n876;
  assign new_n878 = li02 & ~li05;
  assign new_n879 = ~li02 & li05;
  assign new_n880 = ~new_n878 & ~new_n879;
  assign new_n881 = new_n877 & new_n880;
  assign new_n882 = new_n874 & new_n881;
  assign new_n883 = new_n311 & ~new_n882;
  assign li11 = new_n871 | new_n883;
  assign new_n885 = lo12 & ~new_n311;
  assign new_n886 = ~new_n325 & ~new_n360;
  assign new_n887 = ~new_n360 & ~li01;
  assign new_n888 = ~new_n413 & ~new_n887;
  assign new_n889 = new_n325 & ~new_n888;
  assign li29 = new_n886 | new_n889;
  assign new_n891 = lo20 & ~new_n312;
  assign new_n892 = lo20 & ~li00;
  assign new_n893 = ~new_n420 & ~new_n892;
  assign new_n894 = new_n312 & ~new_n893;
  assign li20 = new_n891 | new_n894;
  assign new_n896 = ~li29 & li20;
  assign new_n897 = li29 & ~li20;
  assign new_n898 = ~new_n896 & ~new_n897;
  assign new_n899 = new_n311 & ~new_n898;
  assign li12 = new_n885 | new_n899;
  assign new_n901 = lo13 & ~new_n311;
  assign new_n902 = li00 & ~li01;
  assign new_n903 = ~li00 & li01;
  assign new_n904 = ~new_n902 & ~new_n903;
  assign new_n905 = new_n311 & ~new_n904;
  assign li13 = new_n901 | new_n905;
  assign new_n907 = lo00 & lo15;
  assign new_n908 = lo14 & ~new_n180;
  assign li16 = new_n907 | new_n908;
  assign new_n910 = ~li14 & ~li15;
  assign li18 = lo18 | ~new_n910;
  assign new_n912 = lo18 & new_n311;
  assign po0 = lo16 & new_n912;
  always @ (posedge clock) begin
    lo00 <= li00;
    lo01 <= li01;
    lo02 <= li02;
    lo03 <= li03;
    lo04 <= li04;
    lo05 <= li05;
    lo06 <= li06;
    lo07 <= li07;
    lo08 <= li08;
    lo09 <= li09;
    lo10 <= li10;
    lo11 <= li11;
    lo12 <= li12;
    lo13 <= li13;
    lo14 <= li14;
    lo15 <= li15;
    lo16 <= li16;
    lo17 <= li17;
    lo18 <= li18;
    lo19 <= li19;
    lo20 <= li20;
    lo21 <= li21;
    lo22 <= li22;
    lo23 <= li23;
    lo24 <= li24;
    lo25 <= li25;
    lo26 <= li26;
    lo27 <= li27;
    lo28 <= li28;
    lo29 <= li29;
    lo30 <= li30;
    lo31 <= li31;
    lo32 <= li32;
    lo33 <= li33;
    lo34 <= li34;
    lo35 <= li35;
    lo36 <= li36;
    lo37 <= li37;
    lo38 <= li38;
    lo39 <= li39;
    lo40 <= li40;
    lo41 <= li41;
    lo42 <= li42;
    lo43 <= li43;
    lo44 <= li44;
    lo45 <= li45;
    lo46 <= li46;
    lo47 <= li47;
    lo48 <= li48;
    lo49 <= li49;
    lo50 <= li50;
    lo51 <= li51;
    lo52 <= li52;
    lo53 <= li53;
  end
  initial begin
    lo00 <= 1'b0;
    lo01 <= 1'b0;
    lo02 <= 1'b0;
    lo03 <= 1'b0;
    lo04 <= 1'b0;
    lo05 <= 1'b0;
    lo06 <= 1'b0;
    lo07 <= 1'b0;
    lo08 <= 1'b0;
    lo09 <= 1'b0;
    lo10 <= 1'b0;
    lo11 <= 1'b0;
    lo12 <= 1'b0;
    lo13 <= 1'b0;
    lo14 <= 1'b0;
    lo15 <= 1'b0;
    lo16 <= 1'b0;
    lo17 <= 1'b0;
    lo18 <= 1'b0;
    lo19 <= 1'b0;
    lo20 <= 1'b0;
    lo21 <= 1'b0;
    lo22 <= 1'b0;
    lo23 <= 1'b0;
    lo24 <= 1'b0;
    lo25 <= 1'b0;
    lo26 <= 1'b0;
    lo27 <= 1'b0;
    lo28 <= 1'b0;
    lo29 <= 1'b0;
    lo30 <= 1'b0;
    lo31 <= 1'b0;
    lo32 <= 1'b0;
    lo33 <= 1'b0;
    lo34 <= 1'b0;
    lo35 <= 1'b0;
    lo36 <= 1'b0;
    lo37 <= 1'b0;
    lo38 <= 1'b0;
    lo39 <= 1'b0;
    lo40 <= 1'b0;
    lo41 <= 1'b0;
    lo42 <= 1'b0;
    lo43 <= 1'b0;
    lo44 <= 1'b0;
    lo45 <= 1'b0;
    lo46 <= 1'b0;
    lo47 <= 1'b0;
    lo48 <= 1'b0;
    lo49 <= 1'b0;
    lo50 <= 1'b0;
    lo51 <= 1'b0;
    lo52 <= 1'b0;
    lo53 <= 1'b0;
  end
endmodule


