// Benchmark "multiplier_sc" written by ABC on Fri Jul 19 14:15:06 2024

module multiplier_sc ( clock, 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25,
    po0, po1, po2, po3  );
  input  clock;
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25;
  output po0, po1, po2, po3;
  reg lo00, lo01, lo02, lo03, lo04, lo05, lo06, lo07, lo08, lo09, lo10,
    lo11, lo12, lo13, lo14, lo15, lo16, lo17, lo18, lo19, lo20, lo21, lo22,
    lo23, lo24, lo25, lo26, lo27, lo28, lo29, lo30, lo31, lo32, lo33, lo34,
    lo35, lo36, lo37, lo38, lo39, lo40, lo41, lo42, lo43, lo44, lo45, lo46,
    lo47, lo48, lo49, lo50, lo51, lo52, lo53, lo54, lo55, lo56, lo57, lo58,
    lo59, lo60, lo61, lo62, lo63, lo64, lo65, lo66, lo67, lo68, lo69, lo70,
    lo71, lo72, lo73, lo74, lo75, lo76, lo77, lo78, lo79, lo80, lo81, lo82,
    lo83;
  wire new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n508, new_n509, new_n510, new_n511, new_n512, new_n513, new_n514,
    new_n515, new_n516, new_n517, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1322, new_n1323, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1347, new_n1348, new_n1349, new_n1350, new_n1351,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1359, new_n1360, new_n1361, new_n1362, new_n1363,
    new_n1364, new_n1365, new_n1366, new_n1367, new_n1368, new_n1369,
    new_n1370, new_n1371, new_n1372, new_n1373, new_n1374, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381,
    new_n1382, new_n1383, new_n1384, new_n1385, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422, new_n1423,
    new_n1424, new_n1425, new_n1426, new_n1427, new_n1428, new_n1429,
    new_n1430, new_n1431, new_n1432, new_n1433, new_n1434, new_n1435,
    new_n1436, new_n1437, new_n1438, new_n1439, new_n1440, new_n1441,
    new_n1442, new_n1443, new_n1444, new_n1445, new_n1446, new_n1447,
    new_n1448, new_n1449, new_n1450, new_n1451, new_n1452, new_n1453,
    new_n1454, new_n1455, new_n1456, new_n1457, new_n1458, new_n1459,
    new_n1460, new_n1461, new_n1462, new_n1463, new_n1464, new_n1465,
    new_n1466, new_n1467, new_n1468, new_n1469, new_n1470, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495,
    new_n1496, new_n1497, new_n1498, new_n1499, new_n1500, new_n1501,
    new_n1502, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510, new_n1511, new_n1512, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1720, new_n1721, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727, new_n1728, new_n1729, new_n1730, new_n1731,
    new_n1732, new_n1733, new_n1734, new_n1735, new_n1736, new_n1737,
    new_n1738, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743,
    new_n1744, new_n1745, new_n1746, new_n1747, new_n1748, new_n1749,
    new_n1750, new_n1751, new_n1752, new_n1753, new_n1754, new_n1755,
    new_n1756, new_n1757, new_n1758, new_n1759, new_n1760, new_n1761,
    new_n1762, new_n1763, new_n1764, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1775, new_n1776, new_n1777, new_n1778, new_n1779,
    new_n1780, new_n1781, new_n1782, new_n1783, new_n1784, new_n1785,
    new_n1786, new_n1787, new_n1788, new_n1789, new_n1790, new_n1791,
    new_n1792, new_n1793, new_n1794, new_n1795, new_n1796, new_n1797,
    new_n1798, new_n1800, new_n1801, new_n1802, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1811, new_n1812,
    new_n1813, new_n1814, new_n1815, new_n1816, new_n1817, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1827, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1839,
    new_n1840, new_n1841, new_n1842, new_n1843, new_n1844, new_n1845,
    new_n1846, new_n1847, new_n1848, new_n1849, new_n1850, new_n1852,
    new_n1853, new_n1854, new_n1855, new_n1856, new_n1857, new_n1858,
    new_n1859, new_n1860, new_n1861, new_n1862, new_n1863, new_n1864,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1880, new_n1881, new_n1882, new_n1883, new_n1884,
    new_n1885, new_n1886, new_n1887, new_n1888, new_n1889, new_n1890,
    new_n1891, new_n1892, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906, new_n1907, new_n1909, new_n1910,
    new_n1911, new_n1912, new_n1913, new_n1914, new_n1915, new_n1916,
    new_n1917, new_n1918, new_n1919, new_n1920, new_n1921, new_n1922,
    new_n1923, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1940, new_n1941, new_n1942,
    new_n1943, new_n1944, new_n1945, new_n1946, new_n1947, new_n1948,
    new_n1949, new_n1950, new_n1951, new_n1952, new_n1953, new_n1954,
    new_n1955, new_n1957, new_n1958, new_n1959, new_n1960, new_n1961,
    new_n1962, new_n1963, new_n1964, new_n1965, new_n1966, new_n1967,
    new_n1968, new_n1969, new_n1970, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2003, new_n2004, new_n2005, new_n2006,
    new_n2007, new_n2008, new_n2009, new_n2010, new_n2011, new_n2012,
    new_n2013, new_n2014, new_n2015, new_n2016, new_n2017, new_n2018,
    new_n2019, new_n2020, new_n2021, new_n2022, new_n2023, new_n2024,
    new_n2025, new_n2026, new_n2027, new_n2028, new_n2029, new_n2030,
    new_n2031, new_n2032, new_n2033, new_n2034, new_n2035, new_n2036,
    new_n2037, new_n2038, new_n2039, new_n2040, new_n2041, new_n2042,
    new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049,
    new_n2050, new_n2052, new_n2053, new_n2054, new_n2055, new_n2056,
    new_n2057, new_n2058, new_n2059, new_n2060, new_n2061, new_n2062,
    new_n2063, new_n2064, new_n2065, new_n2067, new_n2068, new_n2069,
    new_n2070, new_n2071, new_n2072, new_n2073, new_n2074, new_n2075,
    new_n2076, new_n2077, new_n2078, new_n2079, new_n2080, new_n2081,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120,
    new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126,
    new_n2127, new_n2128, new_n2130, new_n2131, new_n2132, new_n2133,
    new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139,
    new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2146,
    new_n2147, new_n2148, new_n2149, new_n2150, new_n2151, new_n2152,
    new_n2153, new_n2154, new_n2155, new_n2156, new_n2157, new_n2158,
    new_n2159, new_n2161, new_n2162, new_n2163, new_n2164, new_n2165,
    new_n2166, new_n2167, new_n2168, new_n2169, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190,
    new_n2191, new_n2192, new_n2193, new_n2194, new_n2195, new_n2196,
    new_n2197, new_n2198, new_n2199, new_n2200, new_n2201, new_n2202,
    new_n2203, new_n2204, new_n2205, new_n2206, new_n2207, new_n2208,
    new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214,
    new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220,
    new_n2221, new_n2222, new_n2223, new_n2224, new_n2225, new_n2226,
    new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232,
    new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238,
    new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244,
    new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250,
    new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256,
    new_n2257, new_n2258, new_n2259, new_n2260, new_n2261, new_n2262,
    new_n2263, new_n2264, new_n2265, new_n2266, new_n2267, new_n2268,
    new_n2269, new_n2270, new_n2271, new_n2272, new_n2273, new_n2274,
    new_n2275, new_n2276, new_n2277, new_n2278, new_n2279, new_n2280,
    new_n2281, new_n2282, new_n2283, new_n2284, new_n2285, new_n2286,
    new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304,
    new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316,
    new_n2317, new_n2318, new_n2319, new_n2320, new_n2321, new_n2322,
    new_n2323, new_n2324, new_n2325, new_n2326, new_n2327, new_n2328,
    new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334,
    new_n2335, new_n2336, new_n2337, new_n2338, new_n2339, new_n2340,
    new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2358,
    new_n2359, new_n2360, new_n2361, new_n2362, new_n2363, new_n2364,
    new_n2365, new_n2366, new_n2367, new_n2368, new_n2369, new_n2370,
    new_n2371, new_n2372, new_n2373, new_n2374, new_n2375, new_n2376,
    new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382,
    new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388,
    new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2394,
    new_n2395, new_n2396, new_n2397, new_n2398, new_n2399, new_n2400,
    new_n2401, new_n2402, new_n2403, new_n2404, new_n2405, new_n2406,
    new_n2407, new_n2408, new_n2409, new_n2410, new_n2411, new_n2412,
    new_n2413, new_n2414, new_n2415, new_n2416, new_n2417, new_n2418,
    new_n2419, new_n2420, new_n2421, new_n2422, new_n2423, new_n2424,
    new_n2425, new_n2426, new_n2427, new_n2428, new_n2429, new_n2430,
    new_n2431, new_n2432, new_n2433, new_n2434, new_n2435, new_n2436,
    new_n2437, new_n2438, new_n2439, new_n2440, new_n2441, new_n2442,
    new_n2443, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448,
    new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454,
    new_n2455, new_n2456, new_n2457, new_n2458, new_n2459, new_n2460,
    new_n2461, new_n2462, new_n2463, new_n2464, new_n2465, new_n2466,
    new_n2467, new_n2468, new_n2469, new_n2470, new_n2471, new_n2472,
    new_n2473, new_n2474, new_n2475, new_n2476, new_n2477, new_n2478,
    new_n2479, new_n2480, new_n2481, new_n2482, new_n2483, new_n2484,
    new_n2485, new_n2486, new_n2487, new_n2488, new_n2489, new_n2490,
    new_n2491, new_n2492, new_n2493, new_n2494, new_n2495, new_n2496,
    new_n2497, new_n2498, new_n2499, new_n2500, new_n2501, new_n2502,
    new_n2503, new_n2504, new_n2505, new_n2506, new_n2507, new_n2508,
    new_n2509, new_n2510, new_n2511, new_n2512, new_n2513, new_n2514,
    new_n2515, new_n2516, new_n2517, new_n2518, new_n2519, new_n2520,
    new_n2521, new_n2522, new_n2523, new_n2524, new_n2525, new_n2526,
    new_n2527, new_n2528, new_n2529, new_n2530, new_n2531, new_n2532,
    new_n2533, new_n2534, new_n2535, new_n2536, new_n2537, new_n2538,
    new_n2539, new_n2540, new_n2541, new_n2542, new_n2543, new_n2544,
    new_n2545, new_n2546, new_n2547, new_n2548, new_n2549, new_n2550,
    new_n2551, new_n2552, new_n2553, new_n2554, new_n2555, new_n2556,
    new_n2557, new_n2558, new_n2559, new_n2560, new_n2561, new_n2562,
    new_n2563, new_n2564, new_n2565, new_n2566, new_n2567, new_n2568,
    new_n2569, new_n2570, new_n2571, new_n2572, new_n2573, new_n2574,
    new_n2575, new_n2576, new_n2577, new_n2578, new_n2579, new_n2580,
    new_n2581, new_n2582, new_n2583, new_n2584, new_n2585, new_n2586,
    new_n2587, new_n2588, new_n2589, new_n2590, new_n2591, new_n2592,
    new_n2593, new_n2594, new_n2595, new_n2596, new_n2597, new_n2598,
    new_n2599, new_n2600, new_n2601, new_n2602, new_n2603, new_n2604,
    new_n2605, new_n2606, new_n2607, new_n2608, new_n2609, new_n2610,
    new_n2611, new_n2612, new_n2613, new_n2614, new_n2615, new_n2616,
    new_n2617, new_n2618, new_n2619, new_n2620, new_n2621, new_n2623,
    new_n2624, new_n2625, new_n2626, new_n2627, new_n2628, new_n2629,
    new_n2630, new_n2631, new_n2632, new_n2633, new_n2634, new_n2635,
    new_n2636, new_n2637, new_n2638, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2662, new_n2663, new_n2664, new_n2665, new_n2666, new_n2667,
    new_n2668, new_n2669, new_n2670, new_n2671, new_n2672, new_n2673,
    new_n2674, new_n2675, new_n2676, new_n2677, new_n2679, new_n2680,
    new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686,
    new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692,
    new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698,
    new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2706, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2723, new_n2724,
    new_n2725, new_n2726, new_n2727, new_n2728, new_n2729, new_n2730,
    new_n2731, new_n2732, new_n2733, new_n2734, new_n2735, new_n2736,
    new_n2737, new_n2738, new_n2739, new_n2740, new_n2741, new_n2742,
    new_n2743, new_n2745, new_n2746, new_n2747, new_n2748, new_n2749,
    new_n2750, new_n2751, new_n2752, new_n2753, new_n2754, new_n2755,
    new_n2756, new_n2757, new_n2758, new_n2759, new_n2760, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2790, new_n2791, new_n2792, new_n2793,
    new_n2794, new_n2795, new_n2796, new_n2797, new_n2798, new_n2799,
    new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805,
    new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812,
    new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818,
    new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824,
    new_n2825, new_n2826, new_n2827, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2869,
    new_n2870, new_n2871, new_n2872, new_n2873, new_n2874, new_n2875,
    new_n2876, new_n2877, new_n2878, new_n2879, new_n2880, new_n2881,
    new_n2882, new_n2883, new_n2884, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902, new_n2904, new_n2905, new_n2906, new_n2907,
    new_n2908, new_n2909, new_n2910, new_n2911, new_n2912, new_n2913,
    new_n2914, new_n2915, new_n2916, new_n2917, new_n2918, new_n2919,
    new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926,
    new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932,
    new_n2933, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944, new_n2945,
    new_n2946, new_n2947, new_n2948, new_n2949, new_n2950, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2962, new_n2963, new_n2964, new_n2965,
    new_n2966, new_n2967, new_n2968, new_n2969, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2976, new_n2977, new_n2979, new_n2980,
    new_n2982, new_n2983, new_n2985, new_n2986, new_n2988, new_n2989,
    new_n2991, new_n2992, new_n2994, new_n2995, new_n2997, new_n2998,
    new_n3000, new_n3001, new_n3003, new_n3004, new_n3006, new_n3007,
    new_n3009, new_n3010, new_n3012, new_n3013, new_n3015, new_n3016,
    new_n3018, new_n3019, new_n3021, new_n3022, new_n3024, new_n3025,
    new_n3027, new_n3028, new_n3030, new_n3031, new_n3033, new_n3034,
    new_n3036, new_n3037, new_n3039, new_n3040, new_n3042, new_n3043,
    new_n3045, new_n3046, new_n3048, new_n3049, new_n3051, new_n3052,
    new_n3054, new_n3055, new_n3057, new_n3058, new_n3060, new_n3061,
    new_n3063, new_n3064, new_n3066, new_n3067, new_n3069, new_n3070,
    new_n3072, new_n3073, new_n3075, new_n3077, new_n3079, new_n3081, li00,
    li01, li02, li03, li04, li05, li06, li07, li08, li09, li10, li11, li12,
    li13, li14, li15, li16, li17, li18, li19, li20, li21, li22, li23, li24,
    li25, li26, li27, li28, li29, li30, li31, li32, li33, li34, li35, li36,
    li37, li38, li39, li40, li41, li42, li43, li44, li45, li46, li47, li48,
    li49, li50, li51, li52, li53, li54, li55, li56, li57, li58, li59, li60,
    li61, li62, li63, li64, li65, li66, li67, li68, li69, li70, li71, li72,
    li73, li74, li75, li76, li77, li78, li79, li80, li81, li82, li83;
  assign new_n283 = lo00 & ~lo01;
  assign new_n284 = ~lo00 & lo01;
  assign new_n285 = ~new_n283 & ~new_n284;
  assign new_n286 = ~lo15 & ~new_n285;
  assign new_n287 = ~lo34 & lo43;
  assign new_n288 = lo34 & ~lo43;
  assign new_n289 = ~new_n287 & ~new_n288;
  assign new_n290 = ~lo14 & ~new_n289;
  assign new_n291 = lo05 & ~lo09;
  assign new_n292 = ~lo05 & lo09;
  assign new_n293 = ~new_n291 & ~new_n292;
  assign new_n294 = lo04 & ~lo08;
  assign new_n295 = ~lo04 & lo08;
  assign new_n296 = ~new_n294 & ~new_n295;
  assign new_n297 = new_n293 & new_n296;
  assign new_n298 = lo03 & ~lo07;
  assign new_n299 = ~lo03 & lo07;
  assign new_n300 = ~new_n298 & ~new_n299;
  assign new_n301 = lo02 & ~lo06;
  assign new_n302 = ~lo02 & lo06;
  assign new_n303 = ~new_n301 & ~new_n302;
  assign new_n304 = new_n300 & new_n303;
  assign new_n305 = new_n297 & new_n304;
  assign new_n306 = ~lo13 & ~new_n305;
  assign new_n307 = ~lo12 & lo33;
  assign new_n308 = lo12 & lo75;
  assign new_n309 = ~new_n307 & ~new_n308;
  assign new_n310 = lo33 & new_n309;
  assign new_n311 = ~lo33 & ~new_n309;
  assign new_n312 = ~new_n310 & ~new_n311;
  assign new_n313 = ~lo12 & lo32;
  assign new_n314 = lo12 & lo74;
  assign new_n315 = ~new_n313 & ~new_n314;
  assign new_n316 = lo32 & new_n315;
  assign new_n317 = ~lo32 & ~new_n315;
  assign new_n318 = ~new_n316 & ~new_n317;
  assign new_n319 = new_n312 & new_n318;
  assign new_n320 = ~lo12 & lo31;
  assign new_n321 = lo12 & lo73;
  assign new_n322 = ~new_n320 & ~new_n321;
  assign new_n323 = lo31 & new_n322;
  assign new_n324 = ~lo31 & ~new_n322;
  assign new_n325 = ~new_n323 & ~new_n324;
  assign new_n326 = ~lo12 & lo30;
  assign new_n327 = lo12 & lo72;
  assign new_n328 = ~new_n326 & ~new_n327;
  assign new_n329 = lo30 & new_n328;
  assign new_n330 = ~lo30 & ~new_n328;
  assign new_n331 = ~new_n329 & ~new_n330;
  assign new_n332 = new_n325 & new_n331;
  assign new_n333 = new_n319 & new_n332;
  assign new_n334 = ~lo12 & lo29;
  assign new_n335 = lo12 & lo71;
  assign new_n336 = ~new_n334 & ~new_n335;
  assign new_n337 = lo29 & new_n336;
  assign new_n338 = ~lo29 & ~new_n336;
  assign new_n339 = ~new_n337 & ~new_n338;
  assign new_n340 = ~lo12 & lo28;
  assign new_n341 = lo12 & lo70;
  assign new_n342 = ~new_n340 & ~new_n341;
  assign new_n343 = lo28 & new_n342;
  assign new_n344 = ~lo28 & ~new_n342;
  assign new_n345 = ~new_n343 & ~new_n344;
  assign new_n346 = new_n339 & new_n345;
  assign new_n347 = ~lo12 & lo27;
  assign new_n348 = lo12 & lo69;
  assign new_n349 = ~new_n347 & ~new_n348;
  assign new_n350 = lo27 & new_n349;
  assign new_n351 = ~lo27 & ~new_n349;
  assign new_n352 = ~new_n350 & ~new_n351;
  assign new_n353 = ~lo12 & lo26;
  assign new_n354 = lo12 & lo68;
  assign new_n355 = ~new_n353 & ~new_n354;
  assign new_n356 = lo26 & new_n355;
  assign new_n357 = ~lo26 & ~new_n355;
  assign new_n358 = ~new_n356 & ~new_n357;
  assign new_n359 = new_n352 & new_n358;
  assign new_n360 = new_n346 & new_n359;
  assign new_n361 = new_n333 & new_n360;
  assign new_n362 = ~lo12 & lo25;
  assign new_n363 = lo12 & lo67;
  assign new_n364 = ~new_n362 & ~new_n363;
  assign new_n365 = lo25 & new_n364;
  assign new_n366 = ~lo25 & ~new_n364;
  assign new_n367 = ~new_n365 & ~new_n366;
  assign new_n368 = ~lo12 & lo24;
  assign new_n369 = lo12 & lo66;
  assign new_n370 = ~new_n368 & ~new_n369;
  assign new_n371 = lo24 & new_n370;
  assign new_n372 = ~lo24 & ~new_n370;
  assign new_n373 = ~new_n371 & ~new_n372;
  assign new_n374 = new_n367 & new_n373;
  assign new_n375 = ~lo12 & lo23;
  assign new_n376 = lo12 & lo65;
  assign new_n377 = ~new_n375 & ~new_n376;
  assign new_n378 = lo23 & new_n377;
  assign new_n379 = ~lo23 & ~new_n377;
  assign new_n380 = ~new_n378 & ~new_n379;
  assign new_n381 = ~lo12 & lo22;
  assign new_n382 = lo12 & lo64;
  assign new_n383 = ~new_n381 & ~new_n382;
  assign new_n384 = lo22 & new_n383;
  assign new_n385 = ~lo22 & ~new_n383;
  assign new_n386 = ~new_n384 & ~new_n385;
  assign new_n387 = new_n380 & new_n386;
  assign new_n388 = new_n374 & new_n387;
  assign new_n389 = ~lo12 & lo21;
  assign new_n390 = lo12 & lo63;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = lo21 & new_n391;
  assign new_n393 = ~lo21 & ~new_n391;
  assign new_n394 = ~new_n392 & ~new_n393;
  assign new_n395 = ~lo12 & lo20;
  assign new_n396 = lo12 & lo62;
  assign new_n397 = ~new_n395 & ~new_n396;
  assign new_n398 = lo20 & new_n397;
  assign new_n399 = ~lo20 & ~new_n397;
  assign new_n400 = ~new_n398 & ~new_n399;
  assign new_n401 = new_n394 & new_n400;
  assign new_n402 = ~lo12 & lo19;
  assign new_n403 = lo12 & lo61;
  assign new_n404 = ~new_n402 & ~new_n403;
  assign new_n405 = lo19 & new_n404;
  assign new_n406 = ~lo19 & ~new_n404;
  assign new_n407 = ~new_n405 & ~new_n406;
  assign new_n408 = ~lo12 & lo18;
  assign new_n409 = lo12 & lo60;
  assign new_n410 = ~new_n408 & ~new_n409;
  assign new_n411 = lo18 & new_n410;
  assign new_n412 = ~lo18 & ~new_n410;
  assign new_n413 = ~new_n411 & ~new_n412;
  assign new_n414 = new_n407 & new_n413;
  assign new_n415 = new_n401 & new_n414;
  assign new_n416 = new_n388 & new_n415;
  assign new_n417 = new_n361 & new_n416;
  assign new_n418 = ~lo12 & ~new_n417;
  assign new_n419 = lo42 & ~lo51;
  assign new_n420 = ~lo42 & lo51;
  assign new_n421 = ~new_n419 & ~new_n420;
  assign new_n422 = lo41 & ~lo50;
  assign new_n423 = ~lo41 & lo50;
  assign new_n424 = ~new_n422 & ~new_n423;
  assign new_n425 = new_n421 & new_n424;
  assign new_n426 = lo40 & ~lo49;
  assign new_n427 = ~lo40 & lo49;
  assign new_n428 = ~new_n426 & ~new_n427;
  assign new_n429 = lo39 & ~lo48;
  assign new_n430 = ~lo39 & lo48;
  assign new_n431 = ~new_n429 & ~new_n430;
  assign new_n432 = new_n428 & new_n431;
  assign new_n433 = new_n425 & new_n432;
  assign new_n434 = lo38 & ~lo47;
  assign new_n435 = ~lo38 & lo47;
  assign new_n436 = ~new_n434 & ~new_n435;
  assign new_n437 = lo37 & ~lo46;
  assign new_n438 = ~lo37 & lo46;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign new_n440 = new_n436 & new_n439;
  assign new_n441 = lo36 & ~lo45;
  assign new_n442 = ~lo36 & lo45;
  assign new_n443 = ~new_n441 & ~new_n442;
  assign new_n444 = lo35 & ~lo44;
  assign new_n445 = ~lo35 & lo44;
  assign new_n446 = ~new_n444 & ~new_n445;
  assign new_n447 = new_n443 & new_n446;
  assign new_n448 = new_n440 & new_n447;
  assign new_n449 = new_n433 & new_n448;
  assign new_n450 = ~lo11 & ~new_n449;
  assign new_n451 = ~lo59 & lo83;
  assign new_n452 = lo59 & ~lo83;
  assign new_n453 = ~new_n451 & ~new_n452;
  assign new_n454 = ~lo58 & lo82;
  assign new_n455 = lo58 & ~lo82;
  assign new_n456 = ~new_n454 & ~new_n455;
  assign new_n457 = new_n453 & new_n456;
  assign new_n458 = ~lo57 & lo81;
  assign new_n459 = lo57 & ~lo81;
  assign new_n460 = ~new_n458 & ~new_n459;
  assign new_n461 = ~lo56 & lo80;
  assign new_n462 = lo56 & ~lo80;
  assign new_n463 = ~new_n461 & ~new_n462;
  assign new_n464 = new_n460 & new_n463;
  assign new_n465 = new_n457 & new_n464;
  assign new_n466 = ~lo55 & lo79;
  assign new_n467 = lo55 & ~lo79;
  assign new_n468 = ~new_n466 & ~new_n467;
  assign new_n469 = ~lo54 & lo78;
  assign new_n470 = lo54 & ~lo78;
  assign new_n471 = ~new_n469 & ~new_n470;
  assign new_n472 = new_n468 & new_n471;
  assign new_n473 = ~lo53 & lo77;
  assign new_n474 = lo53 & ~lo77;
  assign new_n475 = ~new_n473 & ~new_n474;
  assign new_n476 = ~lo52 & lo76;
  assign new_n477 = lo52 & ~lo76;
  assign new_n478 = ~new_n476 & ~new_n477;
  assign new_n479 = new_n475 & new_n478;
  assign new_n480 = new_n472 & new_n479;
  assign new_n481 = new_n465 & new_n480;
  assign new_n482 = ~lo10 & ~new_n481;
  assign new_n483 = ~lo17 & ~new_n482;
  assign new_n484 = ~new_n450 & new_n483;
  assign new_n485 = ~new_n418 & new_n484;
  assign new_n486 = ~new_n306 & new_n485;
  assign new_n487 = ~new_n290 & new_n486;
  assign li17 = new_n286 | ~new_n487;
  assign new_n489 = lo51 & lo56;
  assign new_n490 = lo50 & lo57;
  assign new_n491 = lo49 & lo57;
  assign new_n492 = lo48 & lo58;
  assign new_n493 = lo47 & lo59;
  assign new_n494 = ~new_n492 & new_n493;
  assign new_n495 = new_n492 & ~new_n493;
  assign new_n496 = ~new_n494 & ~new_n495;
  assign new_n497 = new_n491 & ~new_n496;
  assign new_n498 = new_n492 & new_n493;
  assign new_n499 = ~new_n497 & ~new_n498;
  assign new_n500 = ~new_n490 & ~new_n499;
  assign new_n501 = new_n490 & new_n499;
  assign new_n502 = ~new_n500 & ~new_n501;
  assign new_n503 = new_n489 & ~new_n502;
  assign new_n504 = new_n490 & ~new_n499;
  assign new_n505 = ~new_n503 & ~new_n504;
  assign new_n506 = ~new_n489 & ~new_n502;
  assign new_n507 = new_n489 & new_n502;
  assign new_n508 = ~new_n506 & ~new_n507;
  assign new_n509 = lo49 & lo58;
  assign new_n510 = lo48 & lo59;
  assign new_n511 = ~new_n509 & new_n510;
  assign new_n512 = new_n509 & ~new_n510;
  assign new_n513 = ~new_n511 & ~new_n512;
  assign new_n514 = ~new_n508 & ~new_n513;
  assign new_n515 = lo51 & lo57;
  assign new_n516 = lo50 & lo58;
  assign new_n517 = new_n509 & new_n510;
  assign new_n518 = ~new_n516 & new_n517;
  assign new_n519 = new_n516 & ~new_n517;
  assign new_n520 = ~new_n518 & ~new_n519;
  assign new_n521 = ~new_n515 & ~new_n520;
  assign new_n522 = new_n515 & new_n520;
  assign new_n523 = ~new_n521 & ~new_n522;
  assign new_n524 = lo49 & lo59;
  assign new_n525 = new_n523 & new_n524;
  assign new_n526 = ~new_n523 & ~new_n524;
  assign new_n527 = ~new_n525 & ~new_n526;
  assign new_n528 = ~new_n514 & ~new_n527;
  assign new_n529 = new_n514 & new_n527;
  assign new_n530 = ~new_n528 & ~new_n529;
  assign new_n531 = ~new_n505 & ~new_n530;
  assign new_n532 = new_n514 & ~new_n527;
  assign new_n533 = ~new_n531 & ~new_n532;
  assign new_n534 = new_n515 & ~new_n520;
  assign new_n535 = new_n516 & new_n517;
  assign new_n536 = ~new_n534 & ~new_n535;
  assign new_n537 = ~new_n523 & new_n524;
  assign new_n538 = lo51 & lo58;
  assign new_n539 = lo50 & lo59;
  assign new_n540 = ~new_n538 & new_n539;
  assign new_n541 = new_n538 & ~new_n539;
  assign new_n542 = ~new_n540 & ~new_n541;
  assign new_n543 = ~new_n537 & ~new_n542;
  assign new_n544 = new_n537 & new_n542;
  assign new_n545 = ~new_n543 & ~new_n544;
  assign new_n546 = new_n536 & ~new_n545;
  assign new_n547 = ~new_n536 & new_n545;
  assign new_n548 = ~new_n546 & ~new_n547;
  assign new_n549 = new_n533 & ~new_n548;
  assign new_n550 = ~new_n533 & new_n548;
  assign new_n551 = ~new_n549 & ~new_n550;
  assign new_n552 = lo51 & lo55;
  assign new_n553 = lo50 & lo56;
  assign new_n554 = lo49 & lo56;
  assign new_n555 = lo48 & lo57;
  assign new_n556 = lo47 & lo58;
  assign new_n557 = ~new_n555 & new_n556;
  assign new_n558 = new_n555 & ~new_n556;
  assign new_n559 = ~new_n557 & ~new_n558;
  assign new_n560 = new_n554 & ~new_n559;
  assign new_n561 = new_n555 & new_n556;
  assign new_n562 = ~new_n560 & ~new_n561;
  assign new_n563 = ~new_n553 & ~new_n562;
  assign new_n564 = new_n553 & new_n562;
  assign new_n565 = ~new_n563 & ~new_n564;
  assign new_n566 = new_n552 & ~new_n565;
  assign new_n567 = new_n553 & ~new_n562;
  assign new_n568 = ~new_n566 & ~new_n567;
  assign new_n569 = ~new_n552 & ~new_n565;
  assign new_n570 = new_n552 & new_n565;
  assign new_n571 = ~new_n569 & ~new_n570;
  assign new_n572 = ~new_n554 & ~new_n559;
  assign new_n573 = new_n554 & new_n559;
  assign new_n574 = ~new_n572 & ~new_n573;
  assign new_n575 = lo46 & lo58;
  assign new_n576 = lo45 & lo59;
  assign new_n577 = new_n575 & new_n576;
  assign new_n578 = lo46 & lo59;
  assign new_n579 = ~new_n577 & new_n578;
  assign new_n580 = new_n577 & ~new_n578;
  assign new_n581 = ~new_n579 & ~new_n580;
  assign new_n582 = ~new_n574 & ~new_n581;
  assign new_n583 = new_n577 & new_n578;
  assign new_n584 = ~new_n582 & ~new_n583;
  assign new_n585 = ~new_n491 & ~new_n496;
  assign new_n586 = new_n491 & new_n496;
  assign new_n587 = ~new_n585 & ~new_n586;
  assign new_n588 = new_n584 & ~new_n587;
  assign new_n589 = ~new_n584 & new_n587;
  assign new_n590 = ~new_n588 & ~new_n589;
  assign new_n591 = ~new_n571 & ~new_n590;
  assign new_n592 = ~new_n584 & ~new_n587;
  assign new_n593 = ~new_n591 & ~new_n592;
  assign new_n594 = new_n508 & ~new_n513;
  assign new_n595 = ~new_n508 & new_n513;
  assign new_n596 = ~new_n594 & ~new_n595;
  assign new_n597 = new_n593 & ~new_n596;
  assign new_n598 = ~new_n593 & new_n596;
  assign new_n599 = ~new_n597 & ~new_n598;
  assign new_n600 = ~new_n568 & ~new_n599;
  assign new_n601 = ~new_n593 & ~new_n596;
  assign new_n602 = ~new_n600 & ~new_n601;
  assign new_n603 = new_n505 & ~new_n530;
  assign new_n604 = ~new_n505 & new_n530;
  assign new_n605 = ~new_n603 & ~new_n604;
  assign new_n606 = new_n602 & ~new_n605;
  assign new_n607 = ~new_n602 & new_n605;
  assign new_n608 = ~new_n606 & ~new_n607;
  assign new_n609 = ~new_n551 & ~new_n608;
  assign new_n610 = lo51 & lo54;
  assign new_n611 = lo50 & lo55;
  assign new_n612 = lo49 & lo55;
  assign new_n613 = lo48 & lo56;
  assign new_n614 = lo47 & lo57;
  assign new_n615 = ~new_n613 & new_n614;
  assign new_n616 = new_n613 & ~new_n614;
  assign new_n617 = ~new_n615 & ~new_n616;
  assign new_n618 = new_n612 & ~new_n617;
  assign new_n619 = new_n613 & new_n614;
  assign new_n620 = ~new_n618 & ~new_n619;
  assign new_n621 = ~new_n611 & ~new_n620;
  assign new_n622 = new_n611 & new_n620;
  assign new_n623 = ~new_n621 & ~new_n622;
  assign new_n624 = new_n610 & ~new_n623;
  assign new_n625 = new_n611 & ~new_n620;
  assign new_n626 = ~new_n624 & ~new_n625;
  assign new_n627 = ~new_n610 & ~new_n623;
  assign new_n628 = new_n610 & new_n623;
  assign new_n629 = ~new_n627 & ~new_n628;
  assign new_n630 = ~new_n612 & ~new_n617;
  assign new_n631 = new_n612 & new_n617;
  assign new_n632 = ~new_n630 & ~new_n631;
  assign new_n633 = lo46 & lo57;
  assign new_n634 = lo45 & lo58;
  assign new_n635 = lo44 & lo59;
  assign new_n636 = ~new_n634 & new_n635;
  assign new_n637 = new_n634 & ~new_n635;
  assign new_n638 = ~new_n636 & ~new_n637;
  assign new_n639 = new_n633 & ~new_n638;
  assign new_n640 = new_n634 & new_n635;
  assign new_n641 = ~new_n639 & ~new_n640;
  assign new_n642 = ~new_n575 & new_n576;
  assign new_n643 = new_n575 & ~new_n576;
  assign new_n644 = ~new_n642 & ~new_n643;
  assign new_n645 = new_n641 & ~new_n644;
  assign new_n646 = ~new_n641 & new_n644;
  assign new_n647 = ~new_n645 & ~new_n646;
  assign new_n648 = ~new_n632 & ~new_n647;
  assign new_n649 = ~new_n641 & ~new_n644;
  assign new_n650 = ~new_n648 & ~new_n649;
  assign new_n651 = new_n574 & ~new_n581;
  assign new_n652 = ~new_n574 & new_n581;
  assign new_n653 = ~new_n651 & ~new_n652;
  assign new_n654 = new_n650 & ~new_n653;
  assign new_n655 = ~new_n650 & new_n653;
  assign new_n656 = ~new_n654 & ~new_n655;
  assign new_n657 = ~new_n629 & ~new_n656;
  assign new_n658 = ~new_n650 & ~new_n653;
  assign new_n659 = ~new_n657 & ~new_n658;
  assign new_n660 = new_n571 & ~new_n590;
  assign new_n661 = ~new_n571 & new_n590;
  assign new_n662 = ~new_n660 & ~new_n661;
  assign new_n663 = new_n659 & ~new_n662;
  assign new_n664 = ~new_n659 & new_n662;
  assign new_n665 = ~new_n663 & ~new_n664;
  assign new_n666 = ~new_n626 & ~new_n665;
  assign new_n667 = ~new_n659 & ~new_n662;
  assign new_n668 = ~new_n666 & ~new_n667;
  assign new_n669 = new_n568 & ~new_n599;
  assign new_n670 = ~new_n568 & new_n599;
  assign new_n671 = ~new_n669 & ~new_n670;
  assign new_n672 = new_n668 & ~new_n671;
  assign new_n673 = ~new_n668 & new_n671;
  assign new_n674 = ~new_n672 & ~new_n673;
  assign new_n675 = lo51 & lo53;
  assign new_n676 = lo50 & lo54;
  assign new_n677 = lo49 & lo54;
  assign new_n678 = lo48 & lo55;
  assign new_n679 = lo47 & lo56;
  assign new_n680 = ~new_n678 & new_n679;
  assign new_n681 = new_n678 & ~new_n679;
  assign new_n682 = ~new_n680 & ~new_n681;
  assign new_n683 = new_n677 & ~new_n682;
  assign new_n684 = new_n678 & new_n679;
  assign new_n685 = ~new_n683 & ~new_n684;
  assign new_n686 = ~new_n676 & ~new_n685;
  assign new_n687 = new_n676 & new_n685;
  assign new_n688 = ~new_n686 & ~new_n687;
  assign new_n689 = new_n675 & ~new_n688;
  assign new_n690 = new_n676 & ~new_n685;
  assign new_n691 = ~new_n689 & ~new_n690;
  assign new_n692 = ~new_n675 & ~new_n688;
  assign new_n693 = new_n675 & new_n688;
  assign new_n694 = ~new_n692 & ~new_n693;
  assign new_n695 = ~new_n677 & ~new_n682;
  assign new_n696 = new_n677 & new_n682;
  assign new_n697 = ~new_n695 & ~new_n696;
  assign new_n698 = lo46 & lo56;
  assign new_n699 = lo45 & lo57;
  assign new_n700 = lo44 & lo58;
  assign new_n701 = ~new_n699 & new_n700;
  assign new_n702 = new_n699 & ~new_n700;
  assign new_n703 = ~new_n701 & ~new_n702;
  assign new_n704 = new_n698 & ~new_n703;
  assign new_n705 = new_n699 & new_n700;
  assign new_n706 = ~new_n704 & ~new_n705;
  assign new_n707 = ~new_n633 & ~new_n638;
  assign new_n708 = new_n633 & new_n638;
  assign new_n709 = ~new_n707 & ~new_n708;
  assign new_n710 = new_n706 & ~new_n709;
  assign new_n711 = ~new_n706 & new_n709;
  assign new_n712 = ~new_n710 & ~new_n711;
  assign new_n713 = ~new_n697 & ~new_n712;
  assign new_n714 = ~new_n706 & ~new_n709;
  assign new_n715 = ~new_n713 & ~new_n714;
  assign new_n716 = new_n632 & ~new_n647;
  assign new_n717 = ~new_n632 & new_n647;
  assign new_n718 = ~new_n716 & ~new_n717;
  assign new_n719 = new_n715 & ~new_n718;
  assign new_n720 = ~new_n715 & new_n718;
  assign new_n721 = ~new_n719 & ~new_n720;
  assign new_n722 = ~new_n694 & ~new_n721;
  assign new_n723 = ~new_n715 & ~new_n718;
  assign new_n724 = ~new_n722 & ~new_n723;
  assign new_n725 = new_n629 & ~new_n656;
  assign new_n726 = ~new_n629 & new_n656;
  assign new_n727 = ~new_n725 & ~new_n726;
  assign new_n728 = new_n724 & ~new_n727;
  assign new_n729 = ~new_n724 & new_n727;
  assign new_n730 = ~new_n728 & ~new_n729;
  assign new_n731 = ~new_n691 & ~new_n730;
  assign new_n732 = ~new_n724 & ~new_n727;
  assign new_n733 = ~new_n731 & ~new_n732;
  assign new_n734 = new_n626 & ~new_n665;
  assign new_n735 = ~new_n626 & new_n665;
  assign new_n736 = ~new_n734 & ~new_n735;
  assign new_n737 = new_n733 & ~new_n736;
  assign new_n738 = ~new_n733 & new_n736;
  assign new_n739 = ~new_n737 & ~new_n738;
  assign new_n740 = ~new_n674 & ~new_n739;
  assign new_n741 = lo51 & lo52;
  assign new_n742 = lo50 & lo53;
  assign new_n743 = lo49 & lo53;
  assign new_n744 = lo48 & lo54;
  assign new_n745 = lo47 & lo55;
  assign new_n746 = ~new_n744 & new_n745;
  assign new_n747 = new_n744 & ~new_n745;
  assign new_n748 = ~new_n746 & ~new_n747;
  assign new_n749 = new_n743 & ~new_n748;
  assign new_n750 = new_n744 & new_n745;
  assign new_n751 = ~new_n749 & ~new_n750;
  assign new_n752 = ~new_n742 & ~new_n751;
  assign new_n753 = new_n742 & new_n751;
  assign new_n754 = ~new_n752 & ~new_n753;
  assign new_n755 = new_n741 & ~new_n754;
  assign new_n756 = new_n742 & ~new_n751;
  assign new_n757 = ~new_n755 & ~new_n756;
  assign new_n758 = ~new_n741 & ~new_n754;
  assign new_n759 = new_n741 & new_n754;
  assign new_n760 = ~new_n758 & ~new_n759;
  assign new_n761 = ~new_n743 & ~new_n748;
  assign new_n762 = new_n743 & new_n748;
  assign new_n763 = ~new_n761 & ~new_n762;
  assign new_n764 = lo46 & lo55;
  assign new_n765 = lo45 & lo56;
  assign new_n766 = lo44 & lo57;
  assign new_n767 = ~new_n765 & new_n766;
  assign new_n768 = new_n765 & ~new_n766;
  assign new_n769 = ~new_n767 & ~new_n768;
  assign new_n770 = new_n764 & ~new_n769;
  assign new_n771 = new_n765 & new_n766;
  assign new_n772 = ~new_n770 & ~new_n771;
  assign new_n773 = ~new_n698 & ~new_n703;
  assign new_n774 = new_n698 & new_n703;
  assign new_n775 = ~new_n773 & ~new_n774;
  assign new_n776 = new_n772 & ~new_n775;
  assign new_n777 = ~new_n772 & new_n775;
  assign new_n778 = ~new_n776 & ~new_n777;
  assign new_n779 = ~new_n763 & ~new_n778;
  assign new_n780 = ~new_n772 & ~new_n775;
  assign new_n781 = ~new_n779 & ~new_n780;
  assign new_n782 = new_n697 & ~new_n712;
  assign new_n783 = ~new_n697 & new_n712;
  assign new_n784 = ~new_n782 & ~new_n783;
  assign new_n785 = new_n781 & ~new_n784;
  assign new_n786 = ~new_n781 & new_n784;
  assign new_n787 = ~new_n785 & ~new_n786;
  assign new_n788 = ~new_n760 & ~new_n787;
  assign new_n789 = ~new_n781 & ~new_n784;
  assign new_n790 = ~new_n788 & ~new_n789;
  assign new_n791 = new_n694 & ~new_n721;
  assign new_n792 = ~new_n694 & new_n721;
  assign new_n793 = ~new_n791 & ~new_n792;
  assign new_n794 = new_n790 & ~new_n793;
  assign new_n795 = ~new_n790 & new_n793;
  assign new_n796 = ~new_n794 & ~new_n795;
  assign new_n797 = ~new_n757 & ~new_n796;
  assign new_n798 = ~new_n790 & ~new_n793;
  assign new_n799 = ~new_n797 & ~new_n798;
  assign new_n800 = new_n691 & ~new_n730;
  assign new_n801 = ~new_n691 & new_n730;
  assign new_n802 = ~new_n800 & ~new_n801;
  assign new_n803 = new_n799 & ~new_n802;
  assign new_n804 = ~new_n799 & new_n802;
  assign new_n805 = ~new_n803 & ~new_n804;
  assign new_n806 = lo50 & lo52;
  assign new_n807 = lo49 & lo52;
  assign new_n808 = lo48 & lo53;
  assign new_n809 = lo47 & lo54;
  assign new_n810 = ~new_n808 & new_n809;
  assign new_n811 = new_n808 & ~new_n809;
  assign new_n812 = ~new_n810 & ~new_n811;
  assign new_n813 = new_n807 & ~new_n812;
  assign new_n814 = new_n808 & new_n809;
  assign new_n815 = ~new_n813 & ~new_n814;
  assign new_n816 = new_n806 & ~new_n815;
  assign new_n817 = ~new_n806 & ~new_n815;
  assign new_n818 = new_n806 & new_n815;
  assign new_n819 = ~new_n817 & ~new_n818;
  assign new_n820 = ~new_n807 & ~new_n812;
  assign new_n821 = new_n807 & new_n812;
  assign new_n822 = ~new_n820 & ~new_n821;
  assign new_n823 = lo46 & lo54;
  assign new_n824 = lo45 & lo55;
  assign new_n825 = lo44 & lo56;
  assign new_n826 = ~new_n824 & new_n825;
  assign new_n827 = new_n824 & ~new_n825;
  assign new_n828 = ~new_n826 & ~new_n827;
  assign new_n829 = new_n823 & ~new_n828;
  assign new_n830 = new_n824 & new_n825;
  assign new_n831 = ~new_n829 & ~new_n830;
  assign new_n832 = ~new_n764 & ~new_n769;
  assign new_n833 = new_n764 & new_n769;
  assign new_n834 = ~new_n832 & ~new_n833;
  assign new_n835 = new_n831 & ~new_n834;
  assign new_n836 = ~new_n831 & new_n834;
  assign new_n837 = ~new_n835 & ~new_n836;
  assign new_n838 = ~new_n822 & ~new_n837;
  assign new_n839 = ~new_n831 & ~new_n834;
  assign new_n840 = ~new_n838 & ~new_n839;
  assign new_n841 = new_n763 & ~new_n778;
  assign new_n842 = ~new_n763 & new_n778;
  assign new_n843 = ~new_n841 & ~new_n842;
  assign new_n844 = new_n840 & ~new_n843;
  assign new_n845 = ~new_n840 & new_n843;
  assign new_n846 = ~new_n844 & ~new_n845;
  assign new_n847 = ~new_n819 & ~new_n846;
  assign new_n848 = ~new_n840 & ~new_n843;
  assign new_n849 = ~new_n847 & ~new_n848;
  assign new_n850 = new_n760 & ~new_n787;
  assign new_n851 = ~new_n760 & new_n787;
  assign new_n852 = ~new_n850 & ~new_n851;
  assign new_n853 = new_n849 & ~new_n852;
  assign new_n854 = ~new_n849 & new_n852;
  assign new_n855 = ~new_n853 & ~new_n854;
  assign new_n856 = new_n816 & ~new_n855;
  assign new_n857 = ~new_n849 & ~new_n852;
  assign new_n858 = ~new_n856 & ~new_n857;
  assign new_n859 = new_n757 & ~new_n796;
  assign new_n860 = ~new_n757 & new_n796;
  assign new_n861 = ~new_n859 & ~new_n860;
  assign new_n862 = new_n858 & ~new_n861;
  assign new_n863 = ~new_n858 & new_n861;
  assign new_n864 = ~new_n862 & ~new_n863;
  assign new_n865 = ~new_n805 & ~new_n864;
  assign new_n866 = new_n740 & new_n865;
  assign new_n867 = lo48 & lo52;
  assign new_n868 = lo47 & lo53;
  assign new_n869 = new_n867 & new_n868;
  assign new_n870 = ~new_n867 & new_n868;
  assign new_n871 = new_n867 & ~new_n868;
  assign new_n872 = ~new_n870 & ~new_n871;
  assign new_n873 = lo46 & lo53;
  assign new_n874 = lo45 & lo54;
  assign new_n875 = lo44 & lo55;
  assign new_n876 = ~new_n874 & new_n875;
  assign new_n877 = new_n874 & ~new_n875;
  assign new_n878 = ~new_n876 & ~new_n877;
  assign new_n879 = new_n873 & ~new_n878;
  assign new_n880 = new_n874 & new_n875;
  assign new_n881 = ~new_n879 & ~new_n880;
  assign new_n882 = ~new_n823 & ~new_n828;
  assign new_n883 = new_n823 & new_n828;
  assign new_n884 = ~new_n882 & ~new_n883;
  assign new_n885 = new_n881 & ~new_n884;
  assign new_n886 = ~new_n881 & new_n884;
  assign new_n887 = ~new_n885 & ~new_n886;
  assign new_n888 = ~new_n872 & ~new_n887;
  assign new_n889 = ~new_n881 & ~new_n884;
  assign new_n890 = ~new_n888 & ~new_n889;
  assign new_n891 = new_n822 & ~new_n837;
  assign new_n892 = ~new_n822 & new_n837;
  assign new_n893 = ~new_n891 & ~new_n892;
  assign new_n894 = new_n890 & ~new_n893;
  assign new_n895 = ~new_n890 & new_n893;
  assign new_n896 = ~new_n894 & ~new_n895;
  assign new_n897 = new_n869 & ~new_n896;
  assign new_n898 = ~new_n890 & ~new_n893;
  assign new_n899 = ~new_n897 & ~new_n898;
  assign new_n900 = new_n819 & ~new_n846;
  assign new_n901 = ~new_n819 & new_n846;
  assign new_n902 = ~new_n900 & ~new_n901;
  assign new_n903 = ~new_n899 & ~new_n902;
  assign new_n904 = ~new_n816 & ~new_n855;
  assign new_n905 = new_n816 & new_n855;
  assign new_n906 = ~new_n904 & ~new_n905;
  assign new_n907 = ~new_n903 & ~new_n906;
  assign new_n908 = new_n903 & new_n906;
  assign new_n909 = ~new_n907 & ~new_n908;
  assign new_n910 = lo47 & lo52;
  assign new_n911 = lo46 & lo52;
  assign new_n912 = lo45 & lo53;
  assign new_n913 = lo44 & lo54;
  assign new_n914 = ~new_n912 & new_n913;
  assign new_n915 = new_n912 & ~new_n913;
  assign new_n916 = ~new_n914 & ~new_n915;
  assign new_n917 = new_n911 & ~new_n916;
  assign new_n918 = new_n912 & new_n913;
  assign new_n919 = ~new_n917 & ~new_n918;
  assign new_n920 = ~new_n873 & ~new_n878;
  assign new_n921 = new_n873 & new_n878;
  assign new_n922 = ~new_n920 & ~new_n921;
  assign new_n923 = new_n919 & ~new_n922;
  assign new_n924 = ~new_n919 & new_n922;
  assign new_n925 = ~new_n923 & ~new_n924;
  assign new_n926 = new_n910 & ~new_n925;
  assign new_n927 = ~new_n919 & ~new_n922;
  assign new_n928 = ~new_n926 & ~new_n927;
  assign new_n929 = new_n872 & ~new_n887;
  assign new_n930 = ~new_n872 & new_n887;
  assign new_n931 = ~new_n929 & ~new_n930;
  assign new_n932 = ~new_n928 & ~new_n931;
  assign new_n933 = ~new_n869 & ~new_n896;
  assign new_n934 = new_n869 & new_n896;
  assign new_n935 = ~new_n933 & ~new_n934;
  assign new_n936 = new_n932 & ~new_n935;
  assign new_n937 = new_n899 & ~new_n902;
  assign new_n938 = ~new_n899 & new_n902;
  assign new_n939 = ~new_n937 & ~new_n938;
  assign new_n940 = ~new_n936 & ~new_n939;
  assign new_n941 = new_n936 & new_n939;
  assign new_n942 = ~new_n940 & ~new_n941;
  assign new_n943 = ~new_n909 & ~new_n942;
  assign new_n944 = lo45 & lo52;
  assign new_n945 = lo44 & lo53;
  assign new_n946 = new_n944 & new_n945;
  assign new_n947 = ~new_n911 & ~new_n916;
  assign new_n948 = new_n911 & new_n916;
  assign new_n949 = ~new_n947 & ~new_n948;
  assign new_n950 = new_n946 & ~new_n949;
  assign new_n951 = ~new_n910 & ~new_n925;
  assign new_n952 = new_n910 & new_n925;
  assign new_n953 = ~new_n951 & ~new_n952;
  assign new_n954 = new_n950 & ~new_n953;
  assign new_n955 = new_n928 & ~new_n931;
  assign new_n956 = ~new_n928 & new_n931;
  assign new_n957 = ~new_n955 & ~new_n956;
  assign new_n958 = new_n954 & ~new_n957;
  assign new_n959 = ~new_n932 & ~new_n935;
  assign new_n960 = new_n932 & new_n935;
  assign new_n961 = ~new_n959 & ~new_n960;
  assign new_n962 = new_n958 & ~new_n961;
  assign new_n963 = new_n943 & new_n962;
  assign new_n964 = new_n936 & ~new_n939;
  assign new_n965 = ~new_n909 & new_n964;
  assign new_n966 = new_n903 & ~new_n906;
  assign new_n967 = ~new_n965 & ~new_n966;
  assign new_n968 = ~new_n963 & new_n967;
  assign new_n969 = new_n866 & ~new_n968;
  assign new_n970 = ~new_n858 & ~new_n861;
  assign new_n971 = ~new_n805 & new_n970;
  assign new_n972 = ~new_n799 & ~new_n802;
  assign new_n973 = ~new_n971 & ~new_n972;
  assign new_n974 = new_n740 & ~new_n973;
  assign new_n975 = ~new_n733 & ~new_n736;
  assign new_n976 = ~new_n674 & new_n975;
  assign new_n977 = ~new_n668 & ~new_n671;
  assign new_n978 = ~new_n976 & ~new_n977;
  assign new_n979 = ~new_n974 & new_n978;
  assign new_n980 = ~new_n969 & new_n979;
  assign new_n981 = new_n609 & ~new_n980;
  assign new_n982 = ~new_n602 & ~new_n605;
  assign new_n983 = ~new_n551 & new_n982;
  assign new_n984 = ~new_n533 & ~new_n548;
  assign new_n985 = ~new_n983 & ~new_n984;
  assign new_n986 = ~new_n981 & new_n985;
  assign new_n987 = ~new_n536 & ~new_n545;
  assign new_n988 = new_n537 & ~new_n542;
  assign new_n989 = ~new_n987 & ~new_n988;
  assign new_n990 = new_n538 & new_n539;
  assign new_n991 = lo51 & lo59;
  assign new_n992 = ~new_n990 & new_n991;
  assign new_n993 = new_n990 & ~new_n991;
  assign new_n994 = ~new_n992 & ~new_n993;
  assign new_n995 = new_n989 & ~new_n994;
  assign new_n996 = ~new_n989 & new_n994;
  assign new_n997 = ~new_n995 & ~new_n996;
  assign new_n998 = ~new_n986 & ~new_n997;
  assign new_n999 = ~new_n989 & ~new_n994;
  assign new_n1000 = ~new_n998 & ~new_n999;
  assign new_n1001 = new_n990 & new_n991;
  assign new_n1002 = new_n1000 & new_n1001;
  assign new_n1003 = ~new_n1000 & ~new_n1001;
  assign new_n1004 = ~new_n1002 & ~new_n1003;
  assign new_n1005 = lo42 & lo80;
  assign new_n1006 = lo41 & lo81;
  assign new_n1007 = lo40 & lo81;
  assign new_n1008 = lo39 & lo82;
  assign new_n1009 = new_n1007 & new_n1008;
  assign new_n1010 = ~new_n1006 & new_n1009;
  assign new_n1011 = new_n1006 & ~new_n1009;
  assign new_n1012 = ~new_n1010 & ~new_n1011;
  assign new_n1013 = new_n1005 & ~new_n1012;
  assign new_n1014 = new_n1006 & new_n1009;
  assign new_n1015 = ~new_n1013 & ~new_n1014;
  assign new_n1016 = ~new_n1005 & ~new_n1012;
  assign new_n1017 = new_n1005 & new_n1012;
  assign new_n1018 = ~new_n1016 & ~new_n1017;
  assign new_n1019 = ~new_n1007 & new_n1008;
  assign new_n1020 = new_n1007 & ~new_n1008;
  assign new_n1021 = ~new_n1019 & ~new_n1020;
  assign new_n1022 = lo38 & lo83;
  assign new_n1023 = ~new_n1021 & new_n1022;
  assign new_n1024 = lo40 & lo82;
  assign new_n1025 = lo39 & lo83;
  assign new_n1026 = ~new_n1024 & new_n1025;
  assign new_n1027 = new_n1024 & ~new_n1025;
  assign new_n1028 = ~new_n1026 & ~new_n1027;
  assign new_n1029 = ~new_n1023 & ~new_n1028;
  assign new_n1030 = new_n1023 & new_n1028;
  assign new_n1031 = ~new_n1029 & ~new_n1030;
  assign new_n1032 = ~new_n1018 & ~new_n1031;
  assign new_n1033 = new_n1023 & ~new_n1028;
  assign new_n1034 = ~new_n1032 & ~new_n1033;
  assign new_n1035 = lo42 & lo81;
  assign new_n1036 = lo41 & lo82;
  assign new_n1037 = new_n1024 & new_n1025;
  assign new_n1038 = ~new_n1036 & new_n1037;
  assign new_n1039 = new_n1036 & ~new_n1037;
  assign new_n1040 = ~new_n1038 & ~new_n1039;
  assign new_n1041 = ~new_n1035 & ~new_n1040;
  assign new_n1042 = new_n1035 & new_n1040;
  assign new_n1043 = ~new_n1041 & ~new_n1042;
  assign new_n1044 = lo40 & lo83;
  assign new_n1045 = new_n1043 & new_n1044;
  assign new_n1046 = ~new_n1043 & ~new_n1044;
  assign new_n1047 = ~new_n1045 & ~new_n1046;
  assign new_n1048 = new_n1034 & ~new_n1047;
  assign new_n1049 = ~new_n1034 & new_n1047;
  assign new_n1050 = ~new_n1048 & ~new_n1049;
  assign new_n1051 = ~new_n1015 & ~new_n1050;
  assign new_n1052 = ~new_n1034 & ~new_n1047;
  assign new_n1053 = ~new_n1051 & ~new_n1052;
  assign new_n1054 = new_n1035 & ~new_n1040;
  assign new_n1055 = new_n1036 & new_n1037;
  assign new_n1056 = ~new_n1054 & ~new_n1055;
  assign new_n1057 = ~new_n1043 & new_n1044;
  assign new_n1058 = lo42 & lo82;
  assign new_n1059 = lo41 & lo83;
  assign new_n1060 = ~new_n1058 & new_n1059;
  assign new_n1061 = new_n1058 & ~new_n1059;
  assign new_n1062 = ~new_n1060 & ~new_n1061;
  assign new_n1063 = ~new_n1057 & ~new_n1062;
  assign new_n1064 = new_n1057 & new_n1062;
  assign new_n1065 = ~new_n1063 & ~new_n1064;
  assign new_n1066 = new_n1056 & ~new_n1065;
  assign new_n1067 = ~new_n1056 & new_n1065;
  assign new_n1068 = ~new_n1066 & ~new_n1067;
  assign new_n1069 = new_n1053 & ~new_n1068;
  assign new_n1070 = ~new_n1053 & new_n1068;
  assign new_n1071 = ~new_n1069 & ~new_n1070;
  assign new_n1072 = lo42 & lo79;
  assign new_n1073 = lo41 & lo80;
  assign new_n1074 = lo40 & lo80;
  assign new_n1075 = lo39 & lo81;
  assign new_n1076 = lo37 & lo83;
  assign new_n1077 = ~new_n1075 & new_n1076;
  assign new_n1078 = new_n1075 & ~new_n1076;
  assign new_n1079 = ~new_n1077 & ~new_n1078;
  assign new_n1080 = new_n1074 & ~new_n1079;
  assign new_n1081 = new_n1075 & new_n1076;
  assign new_n1082 = ~new_n1080 & ~new_n1081;
  assign new_n1083 = ~new_n1073 & ~new_n1082;
  assign new_n1084 = new_n1073 & new_n1082;
  assign new_n1085 = ~new_n1083 & ~new_n1084;
  assign new_n1086 = new_n1072 & ~new_n1085;
  assign new_n1087 = new_n1073 & ~new_n1082;
  assign new_n1088 = ~new_n1086 & ~new_n1087;
  assign new_n1089 = ~new_n1072 & ~new_n1085;
  assign new_n1090 = new_n1072 & new_n1085;
  assign new_n1091 = ~new_n1089 & ~new_n1090;
  assign new_n1092 = ~new_n1074 & ~new_n1079;
  assign new_n1093 = new_n1074 & new_n1079;
  assign new_n1094 = ~new_n1092 & ~new_n1093;
  assign new_n1095 = lo36 & lo83;
  assign new_n1096 = lo38 & lo81;
  assign new_n1097 = new_n1095 & new_n1096;
  assign new_n1098 = lo38 & lo82;
  assign new_n1099 = ~new_n1097 & new_n1098;
  assign new_n1100 = new_n1097 & ~new_n1098;
  assign new_n1101 = ~new_n1099 & ~new_n1100;
  assign new_n1102 = ~new_n1094 & ~new_n1101;
  assign new_n1103 = new_n1097 & new_n1098;
  assign new_n1104 = ~new_n1102 & ~new_n1103;
  assign new_n1105 = new_n1021 & new_n1022;
  assign new_n1106 = ~new_n1021 & ~new_n1022;
  assign new_n1107 = ~new_n1105 & ~new_n1106;
  assign new_n1108 = new_n1104 & ~new_n1107;
  assign new_n1109 = ~new_n1104 & new_n1107;
  assign new_n1110 = ~new_n1108 & ~new_n1109;
  assign new_n1111 = ~new_n1091 & ~new_n1110;
  assign new_n1112 = ~new_n1104 & ~new_n1107;
  assign new_n1113 = ~new_n1111 & ~new_n1112;
  assign new_n1114 = new_n1018 & ~new_n1031;
  assign new_n1115 = ~new_n1018 & new_n1031;
  assign new_n1116 = ~new_n1114 & ~new_n1115;
  assign new_n1117 = new_n1113 & ~new_n1116;
  assign new_n1118 = ~new_n1113 & new_n1116;
  assign new_n1119 = ~new_n1117 & ~new_n1118;
  assign new_n1120 = ~new_n1088 & ~new_n1119;
  assign new_n1121 = ~new_n1113 & ~new_n1116;
  assign new_n1122 = ~new_n1120 & ~new_n1121;
  assign new_n1123 = new_n1015 & ~new_n1050;
  assign new_n1124 = ~new_n1015 & new_n1050;
  assign new_n1125 = ~new_n1123 & ~new_n1124;
  assign new_n1126 = new_n1122 & ~new_n1125;
  assign new_n1127 = ~new_n1122 & new_n1125;
  assign new_n1128 = ~new_n1126 & ~new_n1127;
  assign new_n1129 = ~new_n1071 & ~new_n1128;
  assign new_n1130 = lo42 & lo78;
  assign new_n1131 = lo41 & lo79;
  assign new_n1132 = lo40 & lo79;
  assign new_n1133 = lo39 & lo80;
  assign new_n1134 = lo37 & lo82;
  assign new_n1135 = ~new_n1133 & new_n1134;
  assign new_n1136 = new_n1133 & ~new_n1134;
  assign new_n1137 = ~new_n1135 & ~new_n1136;
  assign new_n1138 = new_n1132 & ~new_n1137;
  assign new_n1139 = new_n1133 & new_n1134;
  assign new_n1140 = ~new_n1138 & ~new_n1139;
  assign new_n1141 = ~new_n1131 & ~new_n1140;
  assign new_n1142 = new_n1131 & new_n1140;
  assign new_n1143 = ~new_n1141 & ~new_n1142;
  assign new_n1144 = new_n1130 & ~new_n1143;
  assign new_n1145 = new_n1131 & ~new_n1140;
  assign new_n1146 = ~new_n1144 & ~new_n1145;
  assign new_n1147 = ~new_n1130 & ~new_n1143;
  assign new_n1148 = new_n1130 & new_n1143;
  assign new_n1149 = ~new_n1147 & ~new_n1148;
  assign new_n1150 = ~new_n1132 & ~new_n1137;
  assign new_n1151 = new_n1132 & new_n1137;
  assign new_n1152 = ~new_n1150 & ~new_n1151;
  assign new_n1153 = lo36 & lo82;
  assign new_n1154 = lo35 & lo83;
  assign new_n1155 = lo38 & lo80;
  assign new_n1156 = ~new_n1154 & new_n1155;
  assign new_n1157 = new_n1154 & ~new_n1155;
  assign new_n1158 = ~new_n1156 & ~new_n1157;
  assign new_n1159 = new_n1153 & ~new_n1158;
  assign new_n1160 = new_n1154 & new_n1155;
  assign new_n1161 = ~new_n1159 & ~new_n1160;
  assign new_n1162 = ~new_n1095 & new_n1096;
  assign new_n1163 = new_n1095 & ~new_n1096;
  assign new_n1164 = ~new_n1162 & ~new_n1163;
  assign new_n1165 = new_n1161 & ~new_n1164;
  assign new_n1166 = ~new_n1161 & new_n1164;
  assign new_n1167 = ~new_n1165 & ~new_n1166;
  assign new_n1168 = ~new_n1152 & ~new_n1167;
  assign new_n1169 = ~new_n1161 & ~new_n1164;
  assign new_n1170 = ~new_n1168 & ~new_n1169;
  assign new_n1171 = new_n1094 & ~new_n1101;
  assign new_n1172 = ~new_n1094 & new_n1101;
  assign new_n1173 = ~new_n1171 & ~new_n1172;
  assign new_n1174 = new_n1170 & ~new_n1173;
  assign new_n1175 = ~new_n1170 & new_n1173;
  assign new_n1176 = ~new_n1174 & ~new_n1175;
  assign new_n1177 = ~new_n1149 & ~new_n1176;
  assign new_n1178 = ~new_n1170 & ~new_n1173;
  assign new_n1179 = ~new_n1177 & ~new_n1178;
  assign new_n1180 = new_n1091 & ~new_n1110;
  assign new_n1181 = ~new_n1091 & new_n1110;
  assign new_n1182 = ~new_n1180 & ~new_n1181;
  assign new_n1183 = new_n1179 & ~new_n1182;
  assign new_n1184 = ~new_n1179 & new_n1182;
  assign new_n1185 = ~new_n1183 & ~new_n1184;
  assign new_n1186 = ~new_n1146 & ~new_n1185;
  assign new_n1187 = ~new_n1179 & ~new_n1182;
  assign new_n1188 = ~new_n1186 & ~new_n1187;
  assign new_n1189 = new_n1088 & ~new_n1119;
  assign new_n1190 = ~new_n1088 & new_n1119;
  assign new_n1191 = ~new_n1189 & ~new_n1190;
  assign new_n1192 = new_n1188 & ~new_n1191;
  assign new_n1193 = ~new_n1188 & new_n1191;
  assign new_n1194 = ~new_n1192 & ~new_n1193;
  assign new_n1195 = lo42 & lo77;
  assign new_n1196 = lo41 & lo78;
  assign new_n1197 = lo40 & lo78;
  assign new_n1198 = lo39 & lo79;
  assign new_n1199 = lo37 & lo81;
  assign new_n1200 = ~new_n1198 & new_n1199;
  assign new_n1201 = new_n1198 & ~new_n1199;
  assign new_n1202 = ~new_n1200 & ~new_n1201;
  assign new_n1203 = new_n1197 & ~new_n1202;
  assign new_n1204 = new_n1198 & new_n1199;
  assign new_n1205 = ~new_n1203 & ~new_n1204;
  assign new_n1206 = ~new_n1196 & ~new_n1205;
  assign new_n1207 = new_n1196 & new_n1205;
  assign new_n1208 = ~new_n1206 & ~new_n1207;
  assign new_n1209 = new_n1195 & ~new_n1208;
  assign new_n1210 = new_n1196 & ~new_n1205;
  assign new_n1211 = ~new_n1209 & ~new_n1210;
  assign new_n1212 = ~new_n1195 & ~new_n1208;
  assign new_n1213 = new_n1195 & new_n1208;
  assign new_n1214 = ~new_n1212 & ~new_n1213;
  assign new_n1215 = ~new_n1197 & ~new_n1202;
  assign new_n1216 = new_n1197 & new_n1202;
  assign new_n1217 = ~new_n1215 & ~new_n1216;
  assign new_n1218 = lo36 & lo81;
  assign new_n1219 = lo35 & lo82;
  assign new_n1220 = lo38 & lo79;
  assign new_n1221 = ~new_n1219 & new_n1220;
  assign new_n1222 = new_n1219 & ~new_n1220;
  assign new_n1223 = ~new_n1221 & ~new_n1222;
  assign new_n1224 = new_n1218 & ~new_n1223;
  assign new_n1225 = new_n1219 & new_n1220;
  assign new_n1226 = ~new_n1224 & ~new_n1225;
  assign new_n1227 = ~new_n1153 & ~new_n1158;
  assign new_n1228 = new_n1153 & new_n1158;
  assign new_n1229 = ~new_n1227 & ~new_n1228;
  assign new_n1230 = new_n1226 & ~new_n1229;
  assign new_n1231 = ~new_n1226 & new_n1229;
  assign new_n1232 = ~new_n1230 & ~new_n1231;
  assign new_n1233 = ~new_n1217 & ~new_n1232;
  assign new_n1234 = ~new_n1226 & ~new_n1229;
  assign new_n1235 = ~new_n1233 & ~new_n1234;
  assign new_n1236 = new_n1152 & ~new_n1167;
  assign new_n1237 = ~new_n1152 & new_n1167;
  assign new_n1238 = ~new_n1236 & ~new_n1237;
  assign new_n1239 = new_n1235 & ~new_n1238;
  assign new_n1240 = ~new_n1235 & new_n1238;
  assign new_n1241 = ~new_n1239 & ~new_n1240;
  assign new_n1242 = ~new_n1214 & ~new_n1241;
  assign new_n1243 = ~new_n1235 & ~new_n1238;
  assign new_n1244 = ~new_n1242 & ~new_n1243;
  assign new_n1245 = new_n1149 & ~new_n1176;
  assign new_n1246 = ~new_n1149 & new_n1176;
  assign new_n1247 = ~new_n1245 & ~new_n1246;
  assign new_n1248 = new_n1244 & ~new_n1247;
  assign new_n1249 = ~new_n1244 & new_n1247;
  assign new_n1250 = ~new_n1248 & ~new_n1249;
  assign new_n1251 = ~new_n1211 & ~new_n1250;
  assign new_n1252 = ~new_n1244 & ~new_n1247;
  assign new_n1253 = ~new_n1251 & ~new_n1252;
  assign new_n1254 = new_n1146 & ~new_n1185;
  assign new_n1255 = ~new_n1146 & new_n1185;
  assign new_n1256 = ~new_n1254 & ~new_n1255;
  assign new_n1257 = new_n1253 & ~new_n1256;
  assign new_n1258 = ~new_n1253 & new_n1256;
  assign new_n1259 = ~new_n1257 & ~new_n1258;
  assign new_n1260 = ~new_n1194 & ~new_n1259;
  assign new_n1261 = lo42 & lo76;
  assign new_n1262 = lo41 & lo77;
  assign new_n1263 = lo40 & lo77;
  assign new_n1264 = lo39 & lo78;
  assign new_n1265 = lo37 & lo80;
  assign new_n1266 = ~new_n1264 & new_n1265;
  assign new_n1267 = new_n1264 & ~new_n1265;
  assign new_n1268 = ~new_n1266 & ~new_n1267;
  assign new_n1269 = new_n1263 & ~new_n1268;
  assign new_n1270 = new_n1264 & new_n1265;
  assign new_n1271 = ~new_n1269 & ~new_n1270;
  assign new_n1272 = ~new_n1262 & ~new_n1271;
  assign new_n1273 = new_n1262 & new_n1271;
  assign new_n1274 = ~new_n1272 & ~new_n1273;
  assign new_n1275 = new_n1261 & ~new_n1274;
  assign new_n1276 = new_n1262 & ~new_n1271;
  assign new_n1277 = ~new_n1275 & ~new_n1276;
  assign new_n1278 = ~new_n1261 & ~new_n1274;
  assign new_n1279 = new_n1261 & new_n1274;
  assign new_n1280 = ~new_n1278 & ~new_n1279;
  assign new_n1281 = ~new_n1263 & ~new_n1268;
  assign new_n1282 = new_n1263 & new_n1268;
  assign new_n1283 = ~new_n1281 & ~new_n1282;
  assign new_n1284 = lo36 & lo80;
  assign new_n1285 = lo35 & lo81;
  assign new_n1286 = lo38 & lo78;
  assign new_n1287 = ~new_n1285 & new_n1286;
  assign new_n1288 = new_n1285 & ~new_n1286;
  assign new_n1289 = ~new_n1287 & ~new_n1288;
  assign new_n1290 = new_n1284 & ~new_n1289;
  assign new_n1291 = new_n1285 & new_n1286;
  assign new_n1292 = ~new_n1290 & ~new_n1291;
  assign new_n1293 = ~new_n1218 & ~new_n1223;
  assign new_n1294 = new_n1218 & new_n1223;
  assign new_n1295 = ~new_n1293 & ~new_n1294;
  assign new_n1296 = new_n1292 & ~new_n1295;
  assign new_n1297 = ~new_n1292 & new_n1295;
  assign new_n1298 = ~new_n1296 & ~new_n1297;
  assign new_n1299 = ~new_n1283 & ~new_n1298;
  assign new_n1300 = ~new_n1292 & ~new_n1295;
  assign new_n1301 = ~new_n1299 & ~new_n1300;
  assign new_n1302 = new_n1217 & ~new_n1232;
  assign new_n1303 = ~new_n1217 & new_n1232;
  assign new_n1304 = ~new_n1302 & ~new_n1303;
  assign new_n1305 = new_n1301 & ~new_n1304;
  assign new_n1306 = ~new_n1301 & new_n1304;
  assign new_n1307 = ~new_n1305 & ~new_n1306;
  assign new_n1308 = ~new_n1280 & ~new_n1307;
  assign new_n1309 = ~new_n1301 & ~new_n1304;
  assign new_n1310 = ~new_n1308 & ~new_n1309;
  assign new_n1311 = new_n1214 & ~new_n1241;
  assign new_n1312 = ~new_n1214 & new_n1241;
  assign new_n1313 = ~new_n1311 & ~new_n1312;
  assign new_n1314 = new_n1310 & ~new_n1313;
  assign new_n1315 = ~new_n1310 & new_n1313;
  assign new_n1316 = ~new_n1314 & ~new_n1315;
  assign new_n1317 = ~new_n1277 & ~new_n1316;
  assign new_n1318 = ~new_n1310 & ~new_n1313;
  assign new_n1319 = ~new_n1317 & ~new_n1318;
  assign new_n1320 = new_n1211 & ~new_n1250;
  assign new_n1321 = ~new_n1211 & new_n1250;
  assign new_n1322 = ~new_n1320 & ~new_n1321;
  assign new_n1323 = new_n1319 & ~new_n1322;
  assign new_n1324 = ~new_n1319 & new_n1322;
  assign new_n1325 = ~new_n1323 & ~new_n1324;
  assign new_n1326 = lo41 & lo76;
  assign new_n1327 = lo40 & lo76;
  assign new_n1328 = lo39 & lo77;
  assign new_n1329 = lo37 & lo79;
  assign new_n1330 = ~new_n1328 & new_n1329;
  assign new_n1331 = new_n1328 & ~new_n1329;
  assign new_n1332 = ~new_n1330 & ~new_n1331;
  assign new_n1333 = new_n1327 & ~new_n1332;
  assign new_n1334 = new_n1328 & new_n1329;
  assign new_n1335 = ~new_n1333 & ~new_n1334;
  assign new_n1336 = new_n1326 & ~new_n1335;
  assign new_n1337 = ~new_n1326 & ~new_n1335;
  assign new_n1338 = new_n1326 & new_n1335;
  assign new_n1339 = ~new_n1337 & ~new_n1338;
  assign new_n1340 = ~new_n1327 & ~new_n1332;
  assign new_n1341 = new_n1327 & new_n1332;
  assign new_n1342 = ~new_n1340 & ~new_n1341;
  assign new_n1343 = lo36 & lo79;
  assign new_n1344 = lo35 & lo80;
  assign new_n1345 = lo38 & lo77;
  assign new_n1346 = ~new_n1344 & new_n1345;
  assign new_n1347 = new_n1344 & ~new_n1345;
  assign new_n1348 = ~new_n1346 & ~new_n1347;
  assign new_n1349 = new_n1343 & ~new_n1348;
  assign new_n1350 = new_n1344 & new_n1345;
  assign new_n1351 = ~new_n1349 & ~new_n1350;
  assign new_n1352 = ~new_n1284 & ~new_n1289;
  assign new_n1353 = new_n1284 & new_n1289;
  assign new_n1354 = ~new_n1352 & ~new_n1353;
  assign new_n1355 = new_n1351 & ~new_n1354;
  assign new_n1356 = ~new_n1351 & new_n1354;
  assign new_n1357 = ~new_n1355 & ~new_n1356;
  assign new_n1358 = ~new_n1342 & ~new_n1357;
  assign new_n1359 = ~new_n1351 & ~new_n1354;
  assign new_n1360 = ~new_n1358 & ~new_n1359;
  assign new_n1361 = new_n1283 & ~new_n1298;
  assign new_n1362 = ~new_n1283 & new_n1298;
  assign new_n1363 = ~new_n1361 & ~new_n1362;
  assign new_n1364 = new_n1360 & ~new_n1363;
  assign new_n1365 = ~new_n1360 & new_n1363;
  assign new_n1366 = ~new_n1364 & ~new_n1365;
  assign new_n1367 = ~new_n1339 & ~new_n1366;
  assign new_n1368 = ~new_n1360 & ~new_n1363;
  assign new_n1369 = ~new_n1367 & ~new_n1368;
  assign new_n1370 = new_n1280 & ~new_n1307;
  assign new_n1371 = ~new_n1280 & new_n1307;
  assign new_n1372 = ~new_n1370 & ~new_n1371;
  assign new_n1373 = new_n1369 & ~new_n1372;
  assign new_n1374 = ~new_n1369 & new_n1372;
  assign new_n1375 = ~new_n1373 & ~new_n1374;
  assign new_n1376 = new_n1336 & ~new_n1375;
  assign new_n1377 = ~new_n1369 & ~new_n1372;
  assign new_n1378 = ~new_n1376 & ~new_n1377;
  assign new_n1379 = new_n1277 & ~new_n1316;
  assign new_n1380 = ~new_n1277 & new_n1316;
  assign new_n1381 = ~new_n1379 & ~new_n1380;
  assign new_n1382 = new_n1378 & ~new_n1381;
  assign new_n1383 = ~new_n1378 & new_n1381;
  assign new_n1384 = ~new_n1382 & ~new_n1383;
  assign new_n1385 = ~new_n1325 & ~new_n1384;
  assign new_n1386 = new_n1260 & new_n1385;
  assign new_n1387 = lo39 & lo76;
  assign new_n1388 = lo37 & lo78;
  assign new_n1389 = new_n1387 & new_n1388;
  assign new_n1390 = ~new_n1387 & new_n1388;
  assign new_n1391 = new_n1387 & ~new_n1388;
  assign new_n1392 = ~new_n1390 & ~new_n1391;
  assign new_n1393 = lo36 & lo78;
  assign new_n1394 = lo35 & lo79;
  assign new_n1395 = lo38 & lo76;
  assign new_n1396 = ~new_n1394 & new_n1395;
  assign new_n1397 = new_n1394 & ~new_n1395;
  assign new_n1398 = ~new_n1396 & ~new_n1397;
  assign new_n1399 = new_n1393 & ~new_n1398;
  assign new_n1400 = new_n1394 & new_n1395;
  assign new_n1401 = ~new_n1399 & ~new_n1400;
  assign new_n1402 = ~new_n1343 & ~new_n1348;
  assign new_n1403 = new_n1343 & new_n1348;
  assign new_n1404 = ~new_n1402 & ~new_n1403;
  assign new_n1405 = new_n1401 & ~new_n1404;
  assign new_n1406 = ~new_n1401 & new_n1404;
  assign new_n1407 = ~new_n1405 & ~new_n1406;
  assign new_n1408 = ~new_n1392 & ~new_n1407;
  assign new_n1409 = ~new_n1401 & ~new_n1404;
  assign new_n1410 = ~new_n1408 & ~new_n1409;
  assign new_n1411 = new_n1342 & ~new_n1357;
  assign new_n1412 = ~new_n1342 & new_n1357;
  assign new_n1413 = ~new_n1411 & ~new_n1412;
  assign new_n1414 = new_n1410 & ~new_n1413;
  assign new_n1415 = ~new_n1410 & new_n1413;
  assign new_n1416 = ~new_n1414 & ~new_n1415;
  assign new_n1417 = new_n1389 & ~new_n1416;
  assign new_n1418 = ~new_n1410 & ~new_n1413;
  assign new_n1419 = ~new_n1417 & ~new_n1418;
  assign new_n1420 = new_n1339 & ~new_n1366;
  assign new_n1421 = ~new_n1339 & new_n1366;
  assign new_n1422 = ~new_n1420 & ~new_n1421;
  assign new_n1423 = ~new_n1419 & ~new_n1422;
  assign new_n1424 = ~new_n1336 & ~new_n1375;
  assign new_n1425 = new_n1336 & new_n1375;
  assign new_n1426 = ~new_n1424 & ~new_n1425;
  assign new_n1427 = ~new_n1423 & ~new_n1426;
  assign new_n1428 = new_n1423 & new_n1426;
  assign new_n1429 = ~new_n1427 & ~new_n1428;
  assign new_n1430 = lo37 & lo77;
  assign new_n1431 = lo36 & lo77;
  assign new_n1432 = lo35 & lo78;
  assign new_n1433 = new_n1431 & new_n1432;
  assign new_n1434 = ~new_n1393 & ~new_n1398;
  assign new_n1435 = new_n1393 & new_n1398;
  assign new_n1436 = ~new_n1434 & ~new_n1435;
  assign new_n1437 = ~new_n1433 & ~new_n1436;
  assign new_n1438 = new_n1433 & new_n1436;
  assign new_n1439 = ~new_n1437 & ~new_n1438;
  assign new_n1440 = new_n1430 & ~new_n1439;
  assign new_n1441 = new_n1433 & ~new_n1436;
  assign new_n1442 = ~new_n1440 & ~new_n1441;
  assign new_n1443 = new_n1392 & ~new_n1407;
  assign new_n1444 = ~new_n1392 & new_n1407;
  assign new_n1445 = ~new_n1443 & ~new_n1444;
  assign new_n1446 = ~new_n1442 & ~new_n1445;
  assign new_n1447 = ~new_n1389 & ~new_n1416;
  assign new_n1448 = new_n1389 & new_n1416;
  assign new_n1449 = ~new_n1447 & ~new_n1448;
  assign new_n1450 = new_n1446 & ~new_n1449;
  assign new_n1451 = new_n1419 & ~new_n1422;
  assign new_n1452 = ~new_n1419 & new_n1422;
  assign new_n1453 = ~new_n1451 & ~new_n1452;
  assign new_n1454 = ~new_n1450 & ~new_n1453;
  assign new_n1455 = new_n1450 & new_n1453;
  assign new_n1456 = ~new_n1454 & ~new_n1455;
  assign new_n1457 = ~new_n1429 & ~new_n1456;
  assign new_n1458 = lo37 & lo76;
  assign new_n1459 = lo36 & lo76;
  assign new_n1460 = lo35 & lo77;
  assign new_n1461 = new_n1459 & new_n1460;
  assign new_n1462 = ~new_n1431 & new_n1432;
  assign new_n1463 = new_n1431 & ~new_n1432;
  assign new_n1464 = ~new_n1462 & ~new_n1463;
  assign new_n1465 = ~new_n1461 & ~new_n1464;
  assign new_n1466 = new_n1461 & new_n1464;
  assign new_n1467 = ~new_n1465 & ~new_n1466;
  assign new_n1468 = new_n1458 & ~new_n1467;
  assign new_n1469 = new_n1461 & ~new_n1464;
  assign new_n1470 = ~new_n1468 & ~new_n1469;
  assign new_n1471 = ~new_n1430 & ~new_n1439;
  assign new_n1472 = new_n1430 & new_n1439;
  assign new_n1473 = ~new_n1471 & ~new_n1472;
  assign new_n1474 = ~new_n1470 & ~new_n1473;
  assign new_n1475 = new_n1442 & ~new_n1445;
  assign new_n1476 = ~new_n1442 & new_n1445;
  assign new_n1477 = ~new_n1475 & ~new_n1476;
  assign new_n1478 = new_n1474 & ~new_n1477;
  assign new_n1479 = ~new_n1446 & ~new_n1449;
  assign new_n1480 = new_n1446 & new_n1449;
  assign new_n1481 = ~new_n1479 & ~new_n1480;
  assign new_n1482 = new_n1478 & ~new_n1481;
  assign new_n1483 = new_n1457 & new_n1482;
  assign new_n1484 = new_n1450 & ~new_n1453;
  assign new_n1485 = ~new_n1429 & new_n1484;
  assign new_n1486 = new_n1423 & ~new_n1426;
  assign new_n1487 = ~new_n1485 & ~new_n1486;
  assign new_n1488 = ~new_n1483 & new_n1487;
  assign new_n1489 = new_n1386 & ~new_n1488;
  assign new_n1490 = ~new_n1378 & ~new_n1381;
  assign new_n1491 = ~new_n1325 & new_n1490;
  assign new_n1492 = ~new_n1319 & ~new_n1322;
  assign new_n1493 = ~new_n1491 & ~new_n1492;
  assign new_n1494 = new_n1260 & ~new_n1493;
  assign new_n1495 = ~new_n1253 & ~new_n1256;
  assign new_n1496 = ~new_n1194 & new_n1495;
  assign new_n1497 = ~new_n1188 & ~new_n1191;
  assign new_n1498 = ~new_n1496 & ~new_n1497;
  assign new_n1499 = ~new_n1494 & new_n1498;
  assign new_n1500 = ~new_n1489 & new_n1499;
  assign new_n1501 = new_n1129 & ~new_n1500;
  assign new_n1502 = ~new_n1122 & ~new_n1125;
  assign new_n1503 = ~new_n1071 & new_n1502;
  assign new_n1504 = ~new_n1053 & ~new_n1068;
  assign new_n1505 = ~new_n1503 & ~new_n1504;
  assign new_n1506 = ~new_n1501 & new_n1505;
  assign new_n1507 = ~new_n1056 & ~new_n1065;
  assign new_n1508 = new_n1057 & ~new_n1062;
  assign new_n1509 = ~new_n1507 & ~new_n1508;
  assign new_n1510 = new_n1058 & new_n1059;
  assign new_n1511 = lo42 & lo83;
  assign new_n1512 = ~new_n1510 & new_n1511;
  assign new_n1513 = new_n1510 & ~new_n1511;
  assign new_n1514 = ~new_n1512 & ~new_n1513;
  assign new_n1515 = new_n1509 & ~new_n1514;
  assign new_n1516 = ~new_n1509 & new_n1514;
  assign new_n1517 = ~new_n1515 & ~new_n1516;
  assign new_n1518 = ~new_n1506 & ~new_n1517;
  assign new_n1519 = ~new_n1509 & ~new_n1514;
  assign new_n1520 = ~new_n1518 & ~new_n1519;
  assign new_n1521 = new_n1510 & new_n1511;
  assign new_n1522 = new_n1520 & new_n1521;
  assign new_n1523 = ~new_n1520 & ~new_n1521;
  assign new_n1524 = ~new_n1522 & ~new_n1523;
  assign new_n1525 = new_n1004 & ~new_n1524;
  assign new_n1526 = ~new_n1004 & new_n1524;
  assign new_n1527 = ~new_n1525 & ~new_n1526;
  assign new_n1528 = new_n986 & ~new_n997;
  assign new_n1529 = ~new_n986 & new_n997;
  assign new_n1530 = ~new_n1528 & ~new_n1529;
  assign new_n1531 = new_n1506 & ~new_n1517;
  assign new_n1532 = ~new_n1506 & new_n1517;
  assign new_n1533 = ~new_n1531 & ~new_n1532;
  assign new_n1534 = new_n1530 & ~new_n1533;
  assign new_n1535 = ~new_n1530 & new_n1533;
  assign new_n1536 = ~new_n1534 & ~new_n1535;
  assign new_n1537 = new_n1527 & new_n1536;
  assign new_n1538 = ~new_n608 & ~new_n980;
  assign new_n1539 = ~new_n982 & ~new_n1538;
  assign new_n1540 = ~new_n551 & new_n1539;
  assign new_n1541 = new_n551 & ~new_n1539;
  assign new_n1542 = ~new_n1540 & ~new_n1541;
  assign new_n1543 = ~new_n1128 & ~new_n1500;
  assign new_n1544 = ~new_n1502 & ~new_n1543;
  assign new_n1545 = ~new_n1071 & new_n1544;
  assign new_n1546 = new_n1071 & ~new_n1544;
  assign new_n1547 = ~new_n1545 & ~new_n1546;
  assign new_n1548 = new_n1542 & ~new_n1547;
  assign new_n1549 = ~new_n1542 & new_n1547;
  assign new_n1550 = ~new_n1548 & ~new_n1549;
  assign new_n1551 = ~new_n608 & new_n980;
  assign new_n1552 = new_n608 & ~new_n980;
  assign new_n1553 = ~new_n1551 & ~new_n1552;
  assign new_n1554 = ~new_n1128 & new_n1500;
  assign new_n1555 = new_n1128 & ~new_n1500;
  assign new_n1556 = ~new_n1554 & ~new_n1555;
  assign new_n1557 = new_n1553 & ~new_n1556;
  assign new_n1558 = ~new_n1553 & new_n1556;
  assign new_n1559 = ~new_n1557 & ~new_n1558;
  assign new_n1560 = new_n1550 & new_n1559;
  assign new_n1561 = new_n1537 & new_n1560;
  assign new_n1562 = new_n865 & ~new_n968;
  assign new_n1563 = new_n973 & ~new_n1562;
  assign new_n1564 = ~new_n739 & ~new_n1563;
  assign new_n1565 = ~new_n975 & ~new_n1564;
  assign new_n1566 = ~new_n674 & new_n1565;
  assign new_n1567 = new_n674 & ~new_n1565;
  assign new_n1568 = ~new_n1566 & ~new_n1567;
  assign new_n1569 = new_n1385 & ~new_n1488;
  assign new_n1570 = new_n1493 & ~new_n1569;
  assign new_n1571 = ~new_n1259 & ~new_n1570;
  assign new_n1572 = ~new_n1495 & ~new_n1571;
  assign new_n1573 = ~new_n1194 & new_n1572;
  assign new_n1574 = new_n1194 & ~new_n1572;
  assign new_n1575 = ~new_n1573 & ~new_n1574;
  assign new_n1576 = new_n1568 & ~new_n1575;
  assign new_n1577 = ~new_n1568 & new_n1575;
  assign new_n1578 = ~new_n1576 & ~new_n1577;
  assign new_n1579 = ~new_n739 & new_n1563;
  assign new_n1580 = new_n739 & ~new_n1563;
  assign new_n1581 = ~new_n1579 & ~new_n1580;
  assign new_n1582 = ~new_n1259 & new_n1570;
  assign new_n1583 = new_n1259 & ~new_n1570;
  assign new_n1584 = ~new_n1582 & ~new_n1583;
  assign new_n1585 = new_n1581 & ~new_n1584;
  assign new_n1586 = ~new_n1581 & new_n1584;
  assign new_n1587 = ~new_n1585 & ~new_n1586;
  assign new_n1588 = new_n1578 & new_n1587;
  assign new_n1589 = ~new_n864 & ~new_n968;
  assign new_n1590 = ~new_n970 & ~new_n1589;
  assign new_n1591 = ~new_n805 & new_n1590;
  assign new_n1592 = new_n805 & ~new_n1590;
  assign new_n1593 = ~new_n1591 & ~new_n1592;
  assign new_n1594 = ~new_n1384 & ~new_n1488;
  assign new_n1595 = ~new_n1490 & ~new_n1594;
  assign new_n1596 = ~new_n1325 & new_n1595;
  assign new_n1597 = new_n1325 & ~new_n1595;
  assign new_n1598 = ~new_n1596 & ~new_n1597;
  assign new_n1599 = new_n1593 & ~new_n1598;
  assign new_n1600 = ~new_n1593 & new_n1598;
  assign new_n1601 = ~new_n1599 & ~new_n1600;
  assign new_n1602 = ~new_n864 & new_n968;
  assign new_n1603 = new_n864 & ~new_n968;
  assign new_n1604 = ~new_n1602 & ~new_n1603;
  assign new_n1605 = ~new_n1384 & new_n1488;
  assign new_n1606 = new_n1384 & ~new_n1488;
  assign new_n1607 = ~new_n1605 & ~new_n1606;
  assign new_n1608 = new_n1604 & ~new_n1607;
  assign new_n1609 = ~new_n1604 & new_n1607;
  assign new_n1610 = ~new_n1608 & ~new_n1609;
  assign new_n1611 = new_n1601 & new_n1610;
  assign new_n1612 = new_n1588 & new_n1611;
  assign new_n1613 = new_n1561 & new_n1612;
  assign new_n1614 = ~new_n942 & new_n962;
  assign new_n1615 = ~new_n964 & ~new_n1614;
  assign new_n1616 = ~new_n909 & new_n1615;
  assign new_n1617 = new_n909 & ~new_n1615;
  assign new_n1618 = ~new_n1616 & ~new_n1617;
  assign new_n1619 = ~new_n1456 & new_n1482;
  assign new_n1620 = ~new_n1484 & ~new_n1619;
  assign new_n1621 = ~new_n1429 & new_n1620;
  assign new_n1622 = new_n1429 & ~new_n1620;
  assign new_n1623 = ~new_n1621 & ~new_n1622;
  assign new_n1624 = new_n1618 & ~new_n1623;
  assign new_n1625 = ~new_n1618 & new_n1623;
  assign new_n1626 = ~new_n1624 & ~new_n1625;
  assign new_n1627 = ~new_n942 & ~new_n962;
  assign new_n1628 = new_n942 & new_n962;
  assign new_n1629 = ~new_n1627 & ~new_n1628;
  assign new_n1630 = ~new_n1456 & ~new_n1482;
  assign new_n1631 = new_n1456 & new_n1482;
  assign new_n1632 = ~new_n1630 & ~new_n1631;
  assign new_n1633 = new_n1629 & ~new_n1632;
  assign new_n1634 = ~new_n1629 & new_n1632;
  assign new_n1635 = ~new_n1633 & ~new_n1634;
  assign new_n1636 = new_n1626 & new_n1635;
  assign new_n1637 = ~new_n958 & ~new_n961;
  assign new_n1638 = new_n958 & new_n961;
  assign new_n1639 = ~new_n1637 & ~new_n1638;
  assign new_n1640 = ~new_n1478 & ~new_n1481;
  assign new_n1641 = new_n1478 & new_n1481;
  assign new_n1642 = ~new_n1640 & ~new_n1641;
  assign new_n1643 = new_n1639 & ~new_n1642;
  assign new_n1644 = ~new_n1639 & new_n1642;
  assign new_n1645 = ~new_n1643 & ~new_n1644;
  assign new_n1646 = ~new_n954 & ~new_n957;
  assign new_n1647 = new_n954 & new_n957;
  assign new_n1648 = ~new_n1646 & ~new_n1647;
  assign new_n1649 = ~new_n1474 & ~new_n1477;
  assign new_n1650 = new_n1474 & new_n1477;
  assign new_n1651 = ~new_n1649 & ~new_n1650;
  assign new_n1652 = new_n1648 & ~new_n1651;
  assign new_n1653 = ~new_n1648 & new_n1651;
  assign new_n1654 = ~new_n1652 & ~new_n1653;
  assign new_n1655 = new_n1645 & new_n1654;
  assign new_n1656 = new_n1636 & new_n1655;
  assign new_n1657 = ~new_n950 & ~new_n953;
  assign new_n1658 = new_n950 & new_n953;
  assign new_n1659 = ~new_n1657 & ~new_n1658;
  assign new_n1660 = new_n1470 & ~new_n1473;
  assign new_n1661 = ~new_n1470 & new_n1473;
  assign new_n1662 = ~new_n1660 & ~new_n1661;
  assign new_n1663 = new_n1659 & ~new_n1662;
  assign new_n1664 = ~new_n1659 & new_n1662;
  assign new_n1665 = ~new_n1663 & ~new_n1664;
  assign new_n1666 = ~new_n946 & ~new_n949;
  assign new_n1667 = new_n946 & new_n949;
  assign new_n1668 = ~new_n1666 & ~new_n1667;
  assign new_n1669 = ~new_n1458 & ~new_n1467;
  assign new_n1670 = new_n1458 & new_n1467;
  assign new_n1671 = ~new_n1669 & ~new_n1670;
  assign new_n1672 = new_n1668 & ~new_n1671;
  assign new_n1673 = ~new_n1668 & new_n1671;
  assign new_n1674 = ~new_n1672 & ~new_n1673;
  assign new_n1675 = new_n1665 & new_n1674;
  assign new_n1676 = ~new_n944 & new_n945;
  assign new_n1677 = new_n944 & ~new_n945;
  assign new_n1678 = ~new_n1676 & ~new_n1677;
  assign new_n1679 = ~new_n1459 & new_n1460;
  assign new_n1680 = new_n1459 & ~new_n1460;
  assign new_n1681 = ~new_n1679 & ~new_n1680;
  assign new_n1682 = new_n1678 & ~new_n1681;
  assign new_n1683 = ~new_n1678 & new_n1681;
  assign new_n1684 = ~new_n1682 & ~new_n1683;
  assign new_n1685 = lo44 & lo52;
  assign new_n1686 = lo35 & lo76;
  assign new_n1687 = ~new_n1685 & new_n1686;
  assign new_n1688 = new_n1685 & ~new_n1686;
  assign new_n1689 = ~new_n1687 & ~new_n1688;
  assign new_n1690 = new_n1684 & new_n1689;
  assign new_n1691 = new_n1675 & new_n1690;
  assign new_n1692 = new_n1656 & new_n1691;
  assign new_n1693 = new_n1613 & new_n1692;
  assign li16 = lo16 | ~new_n1693;
  assign new_n1695 = lo00 & ~lo15;
  assign new_n1696 = lo01 & lo15;
  assign new_n1697 = ~new_n1695 & ~new_n1696;
  assign new_n1698 = lo00 & new_n1697;
  assign new_n1699 = ~li16 & ~new_n1698;
  assign new_n1700 = ~li17 & new_n1699;
  assign new_n1701 = lo00 & ~new_n1700;
  assign new_n1702 = ~lo41 & ~lo42;
  assign new_n1703 = ~lo39 & ~lo40;
  assign new_n1704 = new_n1702 & new_n1703;
  assign new_n1705 = ~lo37 & ~lo38;
  assign new_n1706 = ~lo35 & ~lo36;
  assign new_n1707 = new_n1705 & new_n1706;
  assign new_n1708 = new_n1704 & new_n1707;
  assign new_n1709 = ~lo82 & ~lo83;
  assign new_n1710 = ~lo80 & ~lo81;
  assign new_n1711 = new_n1709 & new_n1710;
  assign new_n1712 = ~lo78 & ~lo79;
  assign new_n1713 = ~lo76 & ~lo77;
  assign new_n1714 = new_n1712 & new_n1713;
  assign new_n1715 = new_n1711 & new_n1714;
  assign new_n1716 = ~new_n1708 & ~new_n1715;
  assign new_n1717 = lo43 & ~new_n1716;
  assign new_n1718 = new_n1700 & new_n1717;
  assign li00 = new_n1701 | new_n1718;
  assign new_n1720 = ~lo10 & ~lo14;
  assign new_n1721 = ~lo11 & new_n1720;
  assign new_n1722 = ~li17 & ~li16;
  assign new_n1723 = ~new_n1721 & new_n1722;
  assign new_n1724 = li00 & ~new_n1723;
  assign new_n1725 = ~lo00 & ~new_n1697;
  assign new_n1726 = ~li16 & ~new_n1725;
  assign new_n1727 = ~li17 & new_n1726;
  assign new_n1728 = ~new_n1697 & ~new_n1727;
  assign new_n1729 = ~lo11 & lo41;
  assign new_n1730 = lo11 & lo50;
  assign new_n1731 = ~new_n1729 & ~new_n1730;
  assign new_n1732 = ~lo11 & lo42;
  assign new_n1733 = lo11 & lo51;
  assign new_n1734 = ~new_n1732 & ~new_n1733;
  assign new_n1735 = new_n1731 & new_n1734;
  assign new_n1736 = ~lo11 & lo39;
  assign new_n1737 = lo11 & lo48;
  assign new_n1738 = ~new_n1736 & ~new_n1737;
  assign new_n1739 = ~lo11 & lo40;
  assign new_n1740 = lo11 & lo49;
  assign new_n1741 = ~new_n1739 & ~new_n1740;
  assign new_n1742 = new_n1738 & new_n1741;
  assign new_n1743 = new_n1735 & new_n1742;
  assign new_n1744 = ~lo11 & lo37;
  assign new_n1745 = lo11 & lo46;
  assign new_n1746 = ~new_n1744 & ~new_n1745;
  assign new_n1747 = ~lo11 & lo38;
  assign new_n1748 = lo11 & lo47;
  assign new_n1749 = ~new_n1747 & ~new_n1748;
  assign new_n1750 = new_n1746 & new_n1749;
  assign new_n1751 = ~lo11 & lo36;
  assign new_n1752 = lo11 & lo45;
  assign new_n1753 = ~new_n1751 & ~new_n1752;
  assign new_n1754 = ~lo11 & lo35;
  assign new_n1755 = lo11 & lo44;
  assign new_n1756 = ~new_n1754 & ~new_n1755;
  assign new_n1757 = new_n1753 & new_n1756;
  assign new_n1758 = new_n1750 & new_n1757;
  assign new_n1759 = new_n1743 & new_n1758;
  assign new_n1760 = ~lo10 & lo82;
  assign new_n1761 = lo10 & lo58;
  assign new_n1762 = ~new_n1760 & ~new_n1761;
  assign new_n1763 = ~lo10 & lo83;
  assign new_n1764 = lo10 & lo59;
  assign new_n1765 = ~new_n1763 & ~new_n1764;
  assign new_n1766 = new_n1762 & new_n1765;
  assign new_n1767 = ~lo10 & lo80;
  assign new_n1768 = lo10 & lo56;
  assign new_n1769 = ~new_n1767 & ~new_n1768;
  assign new_n1770 = ~lo10 & lo81;
  assign new_n1771 = lo10 & lo57;
  assign new_n1772 = ~new_n1770 & ~new_n1771;
  assign new_n1773 = new_n1769 & new_n1772;
  assign new_n1774 = new_n1766 & new_n1773;
  assign new_n1775 = ~lo10 & lo78;
  assign new_n1776 = lo10 & lo54;
  assign new_n1777 = ~new_n1775 & ~new_n1776;
  assign new_n1778 = ~lo10 & lo79;
  assign new_n1779 = lo10 & lo55;
  assign new_n1780 = ~new_n1778 & ~new_n1779;
  assign new_n1781 = new_n1777 & new_n1780;
  assign new_n1782 = ~lo10 & lo76;
  assign new_n1783 = lo10 & lo52;
  assign new_n1784 = ~new_n1782 & ~new_n1783;
  assign new_n1785 = ~lo10 & lo77;
  assign new_n1786 = lo10 & lo53;
  assign new_n1787 = ~new_n1785 & ~new_n1786;
  assign new_n1788 = new_n1784 & new_n1787;
  assign new_n1789 = new_n1781 & new_n1788;
  assign new_n1790 = new_n1774 & new_n1789;
  assign new_n1791 = ~new_n1759 & ~new_n1790;
  assign new_n1792 = ~lo14 & lo43;
  assign new_n1793 = lo14 & lo34;
  assign new_n1794 = ~new_n1792 & ~new_n1793;
  assign new_n1795 = ~new_n1791 & ~new_n1794;
  assign new_n1796 = new_n1727 & new_n1795;
  assign new_n1797 = ~new_n1728 & ~new_n1796;
  assign new_n1798 = new_n1723 & ~new_n1797;
  assign li01 = new_n1724 | new_n1798;
  assign new_n1800 = lo02 & ~new_n1700;
  assign new_n1801 = ~lo02 & lo43;
  assign new_n1802 = new_n1700 & new_n1801;
  assign li02 = new_n1800 | new_n1802;
  assign new_n1804 = lo03 & ~new_n1700;
  assign new_n1805 = ~lo02 & lo03;
  assign new_n1806 = lo02 & ~lo03;
  assign new_n1807 = ~new_n1805 & ~new_n1806;
  assign new_n1808 = lo43 & ~new_n1807;
  assign new_n1809 = new_n1700 & new_n1808;
  assign li03 = new_n1804 | new_n1809;
  assign new_n1811 = lo04 & ~new_n1700;
  assign new_n1812 = lo02 & lo03;
  assign new_n1813 = lo04 & ~new_n1812;
  assign new_n1814 = ~lo04 & new_n1812;
  assign new_n1815 = ~new_n1813 & ~new_n1814;
  assign new_n1816 = lo43 & ~new_n1815;
  assign new_n1817 = new_n1700 & new_n1816;
  assign li04 = new_n1811 | new_n1817;
  assign new_n1819 = lo05 & ~new_n1700;
  assign new_n1820 = lo04 & new_n1812;
  assign new_n1821 = lo05 & ~new_n1820;
  assign new_n1822 = ~lo05 & new_n1820;
  assign new_n1823 = ~new_n1821 & ~new_n1822;
  assign new_n1824 = lo43 & ~new_n1823;
  assign new_n1825 = new_n1700 & new_n1824;
  assign li05 = new_n1819 | new_n1825;
  assign new_n1827 = ~lo13 & ~lo14;
  assign new_n1828 = new_n1722 & ~new_n1827;
  assign new_n1829 = li02 & ~new_n1828;
  assign new_n1830 = lo02 & ~lo13;
  assign new_n1831 = lo06 & lo13;
  assign new_n1832 = ~new_n1830 & ~new_n1831;
  assign new_n1833 = ~new_n1727 & ~new_n1832;
  assign new_n1834 = ~new_n1794 & new_n1832;
  assign new_n1835 = new_n1727 & new_n1834;
  assign new_n1836 = ~new_n1833 & ~new_n1835;
  assign new_n1837 = new_n1828 & ~new_n1836;
  assign li06 = new_n1829 | new_n1837;
  assign new_n1839 = li03 & ~new_n1828;
  assign new_n1840 = lo03 & ~lo13;
  assign new_n1841 = lo07 & lo13;
  assign new_n1842 = ~new_n1840 & ~new_n1841;
  assign new_n1843 = ~new_n1727 & ~new_n1842;
  assign new_n1844 = new_n1832 & ~new_n1842;
  assign new_n1845 = ~new_n1832 & new_n1842;
  assign new_n1846 = ~new_n1844 & ~new_n1845;
  assign new_n1847 = ~new_n1794 & ~new_n1846;
  assign new_n1848 = new_n1727 & new_n1847;
  assign new_n1849 = ~new_n1843 & ~new_n1848;
  assign new_n1850 = new_n1828 & ~new_n1849;
  assign li07 = new_n1839 | new_n1850;
  assign new_n1852 = li04 & ~new_n1828;
  assign new_n1853 = lo04 & ~lo13;
  assign new_n1854 = lo08 & lo13;
  assign new_n1855 = ~new_n1853 & ~new_n1854;
  assign new_n1856 = ~new_n1727 & ~new_n1855;
  assign new_n1857 = ~new_n1832 & ~new_n1842;
  assign new_n1858 = ~new_n1855 & ~new_n1857;
  assign new_n1859 = new_n1855 & new_n1857;
  assign new_n1860 = ~new_n1858 & ~new_n1859;
  assign new_n1861 = ~new_n1794 & ~new_n1860;
  assign new_n1862 = new_n1727 & new_n1861;
  assign new_n1863 = ~new_n1856 & ~new_n1862;
  assign new_n1864 = new_n1828 & ~new_n1863;
  assign li08 = new_n1852 | new_n1864;
  assign new_n1866 = li05 & ~new_n1828;
  assign new_n1867 = lo05 & ~lo13;
  assign new_n1868 = lo09 & lo13;
  assign new_n1869 = ~new_n1867 & ~new_n1868;
  assign new_n1870 = ~new_n1727 & ~new_n1869;
  assign new_n1871 = ~new_n1855 & new_n1857;
  assign new_n1872 = ~new_n1869 & ~new_n1871;
  assign new_n1873 = new_n1869 & new_n1871;
  assign new_n1874 = ~new_n1872 & ~new_n1873;
  assign new_n1875 = ~new_n1794 & ~new_n1874;
  assign new_n1876 = new_n1727 & new_n1875;
  assign new_n1877 = ~new_n1870 & ~new_n1876;
  assign new_n1878 = new_n1828 & ~new_n1877;
  assign li09 = new_n1866 | new_n1878;
  assign new_n1880 = ~new_n1727 & ~new_n1765;
  assign new_n1881 = pi25 & new_n1794;
  assign new_n1882 = pi16 & new_n1881;
  assign new_n1883 = ~new_n1765 & ~new_n1881;
  assign new_n1884 = ~new_n1882 & ~new_n1883;
  assign new_n1885 = new_n1727 & ~new_n1884;
  assign new_n1886 = ~new_n1880 & ~new_n1885;
  assign new_n1887 = lo83 & ~new_n1700;
  assign new_n1888 = pi25 & ~lo43;
  assign new_n1889 = pi08 & new_n1888;
  assign new_n1890 = lo83 & ~new_n1888;
  assign new_n1891 = ~new_n1889 & ~new_n1890;
  assign new_n1892 = new_n1700 & ~new_n1891;
  assign li83 = new_n1887 | new_n1892;
  assign new_n1894 = new_n1886 & li83;
  assign new_n1895 = ~new_n1886 & ~li83;
  assign new_n1896 = ~new_n1894 & ~new_n1895;
  assign new_n1897 = ~new_n1727 & ~new_n1762;
  assign new_n1898 = pi15 & new_n1881;
  assign new_n1899 = ~new_n1762 & ~new_n1881;
  assign new_n1900 = ~new_n1898 & ~new_n1899;
  assign new_n1901 = new_n1727 & ~new_n1900;
  assign new_n1902 = ~new_n1897 & ~new_n1901;
  assign new_n1903 = lo82 & ~new_n1700;
  assign new_n1904 = pi07 & new_n1888;
  assign new_n1905 = lo82 & ~new_n1888;
  assign new_n1906 = ~new_n1904 & ~new_n1905;
  assign new_n1907 = new_n1700 & ~new_n1906;
  assign li82 = new_n1903 | new_n1907;
  assign new_n1909 = new_n1902 & li82;
  assign new_n1910 = ~new_n1902 & ~li82;
  assign new_n1911 = ~new_n1909 & ~new_n1910;
  assign new_n1912 = new_n1896 & new_n1911;
  assign new_n1913 = ~new_n1727 & ~new_n1772;
  assign new_n1914 = pi14 & new_n1881;
  assign new_n1915 = ~new_n1772 & ~new_n1881;
  assign new_n1916 = ~new_n1914 & ~new_n1915;
  assign new_n1917 = new_n1727 & ~new_n1916;
  assign new_n1918 = ~new_n1913 & ~new_n1917;
  assign new_n1919 = lo81 & ~new_n1700;
  assign new_n1920 = pi06 & new_n1888;
  assign new_n1921 = lo81 & ~new_n1888;
  assign new_n1922 = ~new_n1920 & ~new_n1921;
  assign new_n1923 = new_n1700 & ~new_n1922;
  assign li81 = new_n1919 | new_n1923;
  assign new_n1925 = new_n1918 & li81;
  assign new_n1926 = ~new_n1918 & ~li81;
  assign new_n1927 = ~new_n1925 & ~new_n1926;
  assign new_n1928 = ~new_n1727 & ~new_n1769;
  assign new_n1929 = pi13 & new_n1881;
  assign new_n1930 = ~new_n1769 & ~new_n1881;
  assign new_n1931 = ~new_n1929 & ~new_n1930;
  assign new_n1932 = new_n1727 & ~new_n1931;
  assign new_n1933 = ~new_n1928 & ~new_n1932;
  assign new_n1934 = lo80 & ~new_n1700;
  assign new_n1935 = pi05 & new_n1888;
  assign new_n1936 = lo80 & ~new_n1888;
  assign new_n1937 = ~new_n1935 & ~new_n1936;
  assign new_n1938 = new_n1700 & ~new_n1937;
  assign li80 = new_n1934 | new_n1938;
  assign new_n1940 = new_n1933 & li80;
  assign new_n1941 = ~new_n1933 & ~li80;
  assign new_n1942 = ~new_n1940 & ~new_n1941;
  assign new_n1943 = new_n1927 & new_n1942;
  assign new_n1944 = new_n1912 & new_n1943;
  assign new_n1945 = ~new_n1727 & ~new_n1780;
  assign new_n1946 = pi12 & new_n1881;
  assign new_n1947 = ~new_n1780 & ~new_n1881;
  assign new_n1948 = ~new_n1946 & ~new_n1947;
  assign new_n1949 = new_n1727 & ~new_n1948;
  assign new_n1950 = ~new_n1945 & ~new_n1949;
  assign new_n1951 = lo79 & ~new_n1700;
  assign new_n1952 = pi04 & new_n1888;
  assign new_n1953 = lo79 & ~new_n1888;
  assign new_n1954 = ~new_n1952 & ~new_n1953;
  assign new_n1955 = new_n1700 & ~new_n1954;
  assign li79 = new_n1951 | new_n1955;
  assign new_n1957 = new_n1950 & li79;
  assign new_n1958 = ~new_n1950 & ~li79;
  assign new_n1959 = ~new_n1957 & ~new_n1958;
  assign new_n1960 = ~new_n1727 & ~new_n1777;
  assign new_n1961 = pi11 & new_n1881;
  assign new_n1962 = ~new_n1777 & ~new_n1881;
  assign new_n1963 = ~new_n1961 & ~new_n1962;
  assign new_n1964 = new_n1727 & ~new_n1963;
  assign new_n1965 = ~new_n1960 & ~new_n1964;
  assign new_n1966 = lo78 & ~new_n1700;
  assign new_n1967 = pi03 & new_n1888;
  assign new_n1968 = lo78 & ~new_n1888;
  assign new_n1969 = ~new_n1967 & ~new_n1968;
  assign new_n1970 = new_n1700 & ~new_n1969;
  assign li78 = new_n1966 | new_n1970;
  assign new_n1972 = new_n1965 & li78;
  assign new_n1973 = ~new_n1965 & ~li78;
  assign new_n1974 = ~new_n1972 & ~new_n1973;
  assign new_n1975 = new_n1959 & new_n1974;
  assign new_n1976 = ~new_n1727 & ~new_n1787;
  assign new_n1977 = pi10 & new_n1881;
  assign new_n1978 = ~new_n1787 & ~new_n1881;
  assign new_n1979 = ~new_n1977 & ~new_n1978;
  assign new_n1980 = new_n1727 & ~new_n1979;
  assign new_n1981 = ~new_n1976 & ~new_n1980;
  assign new_n1982 = lo77 & ~new_n1700;
  assign new_n1983 = pi02 & new_n1888;
  assign new_n1984 = lo77 & ~new_n1888;
  assign new_n1985 = ~new_n1983 & ~new_n1984;
  assign new_n1986 = new_n1700 & ~new_n1985;
  assign li77 = new_n1982 | new_n1986;
  assign new_n1988 = new_n1981 & li77;
  assign new_n1989 = ~new_n1981 & ~li77;
  assign new_n1990 = ~new_n1988 & ~new_n1989;
  assign new_n1991 = ~new_n1727 & ~new_n1784;
  assign new_n1992 = pi09 & new_n1881;
  assign new_n1993 = ~new_n1784 & ~new_n1881;
  assign new_n1994 = ~new_n1992 & ~new_n1993;
  assign new_n1995 = new_n1727 & ~new_n1994;
  assign new_n1996 = ~new_n1991 & ~new_n1995;
  assign new_n1997 = lo76 & ~new_n1700;
  assign new_n1998 = pi01 & new_n1888;
  assign new_n1999 = lo76 & ~new_n1888;
  assign new_n2000 = ~new_n1998 & ~new_n1999;
  assign new_n2001 = new_n1700 & ~new_n2000;
  assign li76 = new_n1997 | new_n2001;
  assign new_n2003 = new_n1996 & li76;
  assign new_n2004 = ~new_n1996 & ~li76;
  assign new_n2005 = ~new_n2003 & ~new_n2004;
  assign new_n2006 = new_n1990 & new_n2005;
  assign new_n2007 = new_n1975 & new_n2006;
  assign new_n2008 = new_n1944 & new_n2007;
  assign new_n2009 = pi08 & ~pi16;
  assign new_n2010 = ~pi08 & pi16;
  assign new_n2011 = ~new_n2009 & ~new_n2010;
  assign new_n2012 = pi07 & ~pi15;
  assign new_n2013 = ~pi07 & pi15;
  assign new_n2014 = ~new_n2012 & ~new_n2013;
  assign new_n2015 = new_n2011 & new_n2014;
  assign new_n2016 = pi06 & ~pi14;
  assign new_n2017 = ~pi06 & pi14;
  assign new_n2018 = ~new_n2016 & ~new_n2017;
  assign new_n2019 = pi05 & ~pi13;
  assign new_n2020 = ~pi05 & pi13;
  assign new_n2021 = ~new_n2019 & ~new_n2020;
  assign new_n2022 = new_n2018 & new_n2021;
  assign new_n2023 = new_n2015 & new_n2022;
  assign new_n2024 = pi04 & ~pi12;
  assign new_n2025 = ~pi04 & pi12;
  assign new_n2026 = ~new_n2024 & ~new_n2025;
  assign new_n2027 = pi03 & ~pi11;
  assign new_n2028 = ~pi03 & pi11;
  assign new_n2029 = ~new_n2027 & ~new_n2028;
  assign new_n2030 = new_n2026 & new_n2029;
  assign new_n2031 = pi02 & ~pi10;
  assign new_n2032 = ~pi02 & pi10;
  assign new_n2033 = ~new_n2031 & ~new_n2032;
  assign new_n2034 = pi01 & ~pi09;
  assign new_n2035 = ~pi01 & pi09;
  assign new_n2036 = ~new_n2034 & ~new_n2035;
  assign new_n2037 = new_n2033 & new_n2036;
  assign new_n2038 = new_n2030 & new_n2037;
  assign new_n2039 = new_n2023 & new_n2038;
  assign new_n2040 = new_n1720 & new_n2039;
  assign new_n2041 = new_n1722 & ~new_n2040;
  assign new_n2042 = ~new_n2008 & new_n2041;
  assign li10 = new_n1700 & new_n2042;
  assign new_n2044 = ~new_n1727 & ~new_n1734;
  assign new_n2045 = pi24 & new_n1881;
  assign new_n2046 = new_n1727 & new_n2045;
  assign new_n2047 = ~new_n2044 & ~new_n2046;
  assign new_n2048 = lo42 & ~new_n1700;
  assign new_n2049 = pi24 & new_n1888;
  assign new_n2050 = new_n1700 & new_n2049;
  assign li42 = new_n2048 | new_n2050;
  assign new_n2052 = new_n2047 & li42;
  assign new_n2053 = ~new_n2047 & ~li42;
  assign new_n2054 = ~new_n2052 & ~new_n2053;
  assign new_n2055 = ~new_n1727 & ~new_n1731;
  assign new_n2056 = pi23 & new_n1881;
  assign new_n2057 = ~new_n1734 & ~new_n1881;
  assign new_n2058 = ~new_n2056 & ~new_n2057;
  assign new_n2059 = new_n1727 & ~new_n2058;
  assign new_n2060 = ~new_n2055 & ~new_n2059;
  assign new_n2061 = lo41 & ~new_n1700;
  assign new_n2062 = pi23 & new_n1888;
  assign new_n2063 = lo42 & ~new_n1888;
  assign new_n2064 = ~new_n2062 & ~new_n2063;
  assign new_n2065 = new_n1700 & ~new_n2064;
  assign li41 = new_n2061 | new_n2065;
  assign new_n2067 = new_n2060 & li41;
  assign new_n2068 = ~new_n2060 & ~li41;
  assign new_n2069 = ~new_n2067 & ~new_n2068;
  assign new_n2070 = new_n2054 & new_n2069;
  assign new_n2071 = ~new_n1727 & ~new_n1741;
  assign new_n2072 = pi22 & new_n1881;
  assign new_n2073 = ~new_n1731 & ~new_n1881;
  assign new_n2074 = ~new_n2072 & ~new_n2073;
  assign new_n2075 = new_n1727 & ~new_n2074;
  assign new_n2076 = ~new_n2071 & ~new_n2075;
  assign new_n2077 = lo40 & ~new_n1700;
  assign new_n2078 = pi22 & new_n1888;
  assign new_n2079 = lo41 & ~new_n1888;
  assign new_n2080 = ~new_n2078 & ~new_n2079;
  assign new_n2081 = new_n1700 & ~new_n2080;
  assign li40 = new_n2077 | new_n2081;
  assign new_n2083 = new_n2076 & li40;
  assign new_n2084 = ~new_n2076 & ~li40;
  assign new_n2085 = ~new_n2083 & ~new_n2084;
  assign new_n2086 = ~new_n1727 & ~new_n1738;
  assign new_n2087 = pi21 & new_n1881;
  assign new_n2088 = ~new_n1741 & ~new_n1881;
  assign new_n2089 = ~new_n2087 & ~new_n2088;
  assign new_n2090 = new_n1727 & ~new_n2089;
  assign new_n2091 = ~new_n2086 & ~new_n2090;
  assign new_n2092 = lo39 & ~new_n1700;
  assign new_n2093 = pi21 & new_n1888;
  assign new_n2094 = lo40 & ~new_n1888;
  assign new_n2095 = ~new_n2093 & ~new_n2094;
  assign new_n2096 = new_n1700 & ~new_n2095;
  assign li39 = new_n2092 | new_n2096;
  assign new_n2098 = new_n2091 & li39;
  assign new_n2099 = ~new_n2091 & ~li39;
  assign new_n2100 = ~new_n2098 & ~new_n2099;
  assign new_n2101 = new_n2085 & new_n2100;
  assign new_n2102 = new_n2070 & new_n2101;
  assign new_n2103 = ~new_n1727 & ~new_n1749;
  assign new_n2104 = pi20 & new_n1881;
  assign new_n2105 = ~new_n1738 & ~new_n1881;
  assign new_n2106 = ~new_n2104 & ~new_n2105;
  assign new_n2107 = new_n1727 & ~new_n2106;
  assign new_n2108 = ~new_n2103 & ~new_n2107;
  assign new_n2109 = lo38 & ~new_n1700;
  assign new_n2110 = pi20 & new_n1888;
  assign new_n2111 = lo39 & ~new_n1888;
  assign new_n2112 = ~new_n2110 & ~new_n2111;
  assign new_n2113 = new_n1700 & ~new_n2112;
  assign li38 = new_n2109 | new_n2113;
  assign new_n2115 = new_n2108 & li38;
  assign new_n2116 = ~new_n2108 & ~li38;
  assign new_n2117 = ~new_n2115 & ~new_n2116;
  assign new_n2118 = ~new_n1727 & ~new_n1746;
  assign new_n2119 = pi19 & new_n1881;
  assign new_n2120 = ~new_n1749 & ~new_n1881;
  assign new_n2121 = ~new_n2119 & ~new_n2120;
  assign new_n2122 = new_n1727 & ~new_n2121;
  assign new_n2123 = ~new_n2118 & ~new_n2122;
  assign new_n2124 = lo37 & ~new_n1700;
  assign new_n2125 = pi19 & new_n1888;
  assign new_n2126 = lo38 & ~new_n1888;
  assign new_n2127 = ~new_n2125 & ~new_n2126;
  assign new_n2128 = new_n1700 & ~new_n2127;
  assign li37 = new_n2124 | new_n2128;
  assign new_n2130 = new_n2123 & li37;
  assign new_n2131 = ~new_n2123 & ~li37;
  assign new_n2132 = ~new_n2130 & ~new_n2131;
  assign new_n2133 = new_n2117 & new_n2132;
  assign new_n2134 = ~new_n1727 & ~new_n1753;
  assign new_n2135 = pi18 & new_n1881;
  assign new_n2136 = ~new_n1746 & ~new_n1881;
  assign new_n2137 = ~new_n2135 & ~new_n2136;
  assign new_n2138 = new_n1727 & ~new_n2137;
  assign new_n2139 = ~new_n2134 & ~new_n2138;
  assign new_n2140 = lo36 & ~new_n1700;
  assign new_n2141 = pi18 & new_n1888;
  assign new_n2142 = lo37 & ~new_n1888;
  assign new_n2143 = ~new_n2141 & ~new_n2142;
  assign new_n2144 = new_n1700 & ~new_n2143;
  assign li36 = new_n2140 | new_n2144;
  assign new_n2146 = new_n2139 & li36;
  assign new_n2147 = ~new_n2139 & ~li36;
  assign new_n2148 = ~new_n2146 & ~new_n2147;
  assign new_n2149 = ~new_n1727 & ~new_n1756;
  assign new_n2150 = pi17 & new_n1881;
  assign new_n2151 = ~new_n1753 & ~new_n1881;
  assign new_n2152 = ~new_n2150 & ~new_n2151;
  assign new_n2153 = new_n1727 & ~new_n2152;
  assign new_n2154 = ~new_n2149 & ~new_n2153;
  assign new_n2155 = lo35 & ~new_n1700;
  assign new_n2156 = pi17 & new_n1888;
  assign new_n2157 = lo36 & ~new_n1888;
  assign new_n2158 = ~new_n2156 & ~new_n2157;
  assign new_n2159 = new_n1700 & ~new_n2158;
  assign li35 = new_n2155 | new_n2159;
  assign new_n2161 = new_n2154 & li35;
  assign new_n2162 = ~new_n2154 & ~li35;
  assign new_n2163 = ~new_n2161 & ~new_n2162;
  assign new_n2164 = new_n2148 & new_n2163;
  assign new_n2165 = new_n2133 & new_n2164;
  assign new_n2166 = new_n2102 & new_n2165;
  assign new_n2167 = ~lo11 & ~lo14;
  assign new_n2168 = new_n1722 & ~new_n2167;
  assign new_n2169 = ~new_n2166 & new_n2168;
  assign li11 = new_n1700 & new_n2169;
  assign new_n2171 = ~new_n309 & ~new_n1727;
  assign new_n2172 = ~new_n1784 & new_n1832;
  assign new_n2173 = new_n1842 & new_n2172;
  assign new_n2174 = new_n1855 & new_n2173;
  assign new_n2175 = new_n1869 & new_n2174;
  assign new_n2176 = ~new_n1756 & new_n2175;
  assign new_n2177 = ~new_n410 & new_n2176;
  assign new_n2178 = ~new_n1784 & ~new_n1832;
  assign new_n2179 = ~new_n1787 & new_n1832;
  assign new_n2180 = ~new_n2178 & ~new_n2179;
  assign new_n2181 = new_n1842 & ~new_n2180;
  assign new_n2182 = new_n1855 & new_n2181;
  assign new_n2183 = new_n1869 & new_n2182;
  assign new_n2184 = ~new_n1756 & new_n2183;
  assign new_n2185 = new_n404 & new_n2184;
  assign new_n2186 = ~new_n404 & ~new_n2184;
  assign new_n2187 = ~new_n2185 & ~new_n2186;
  assign new_n2188 = new_n2177 & ~new_n2187;
  assign new_n2189 = ~new_n404 & new_n2184;
  assign new_n2190 = ~new_n2188 & ~new_n2189;
  assign new_n2191 = ~new_n1842 & new_n2172;
  assign new_n2192 = ~new_n1787 & ~new_n1832;
  assign new_n2193 = ~new_n1777 & new_n1832;
  assign new_n2194 = ~new_n2192 & ~new_n2193;
  assign new_n2195 = new_n1842 & ~new_n2194;
  assign new_n2196 = ~new_n2191 & ~new_n2195;
  assign new_n2197 = new_n1855 & ~new_n2196;
  assign new_n2198 = new_n1869 & new_n2197;
  assign new_n2199 = ~new_n1756 & new_n2198;
  assign new_n2200 = new_n397 & new_n2199;
  assign new_n2201 = ~new_n397 & ~new_n2199;
  assign new_n2202 = ~new_n2200 & ~new_n2201;
  assign new_n2203 = ~new_n1842 & ~new_n2180;
  assign new_n2204 = ~new_n1777 & ~new_n1832;
  assign new_n2205 = ~new_n1780 & new_n1832;
  assign new_n2206 = ~new_n2204 & ~new_n2205;
  assign new_n2207 = new_n1842 & ~new_n2206;
  assign new_n2208 = ~new_n2203 & ~new_n2207;
  assign new_n2209 = new_n1855 & ~new_n2208;
  assign new_n2210 = new_n1869 & new_n2209;
  assign new_n2211 = ~new_n1756 & new_n2210;
  assign new_n2212 = new_n391 & new_n2211;
  assign new_n2213 = ~new_n391 & ~new_n2211;
  assign new_n2214 = ~new_n2212 & ~new_n2213;
  assign new_n2215 = ~new_n2202 & ~new_n2214;
  assign new_n2216 = ~new_n2190 & new_n2215;
  assign new_n2217 = ~new_n397 & new_n2199;
  assign new_n2218 = ~new_n2214 & new_n2217;
  assign new_n2219 = ~new_n391 & new_n2211;
  assign new_n2220 = ~new_n2218 & ~new_n2219;
  assign new_n2221 = ~new_n2216 & new_n2220;
  assign new_n2222 = ~new_n1855 & new_n2173;
  assign new_n2223 = ~new_n1842 & ~new_n2194;
  assign new_n2224 = ~new_n1780 & ~new_n1832;
  assign new_n2225 = ~new_n1769 & new_n1832;
  assign new_n2226 = ~new_n2224 & ~new_n2225;
  assign new_n2227 = new_n1842 & ~new_n2226;
  assign new_n2228 = ~new_n2223 & ~new_n2227;
  assign new_n2229 = new_n1855 & ~new_n2228;
  assign new_n2230 = ~new_n2222 & ~new_n2229;
  assign new_n2231 = new_n1869 & ~new_n2230;
  assign new_n2232 = ~new_n1756 & new_n2231;
  assign new_n2233 = new_n383 & new_n2232;
  assign new_n2234 = ~new_n383 & ~new_n2232;
  assign new_n2235 = ~new_n2233 & ~new_n2234;
  assign new_n2236 = ~new_n1855 & new_n2181;
  assign new_n2237 = ~new_n1842 & ~new_n2206;
  assign new_n2238 = ~new_n1769 & ~new_n1832;
  assign new_n2239 = ~new_n1772 & new_n1832;
  assign new_n2240 = ~new_n2238 & ~new_n2239;
  assign new_n2241 = new_n1842 & ~new_n2240;
  assign new_n2242 = ~new_n2237 & ~new_n2241;
  assign new_n2243 = new_n1855 & ~new_n2242;
  assign new_n2244 = ~new_n2236 & ~new_n2243;
  assign new_n2245 = new_n1869 & ~new_n2244;
  assign new_n2246 = ~new_n1756 & new_n2245;
  assign new_n2247 = new_n377 & new_n2246;
  assign new_n2248 = ~new_n377 & ~new_n2246;
  assign new_n2249 = ~new_n2247 & ~new_n2248;
  assign new_n2250 = ~new_n2235 & ~new_n2249;
  assign new_n2251 = ~new_n1855 & ~new_n2196;
  assign new_n2252 = ~new_n1842 & ~new_n2226;
  assign new_n2253 = ~new_n1772 & ~new_n1832;
  assign new_n2254 = ~new_n1762 & new_n1832;
  assign new_n2255 = ~new_n2253 & ~new_n2254;
  assign new_n2256 = new_n1842 & ~new_n2255;
  assign new_n2257 = ~new_n2252 & ~new_n2256;
  assign new_n2258 = new_n1855 & ~new_n2257;
  assign new_n2259 = ~new_n2251 & ~new_n2258;
  assign new_n2260 = new_n1869 & ~new_n2259;
  assign new_n2261 = ~new_n1756 & new_n2260;
  assign new_n2262 = new_n370 & new_n2261;
  assign new_n2263 = ~new_n370 & ~new_n2261;
  assign new_n2264 = ~new_n2262 & ~new_n2263;
  assign new_n2265 = ~new_n1855 & ~new_n2208;
  assign new_n2266 = ~new_n1842 & ~new_n2240;
  assign new_n2267 = ~new_n1762 & ~new_n1832;
  assign new_n2268 = ~new_n1765 & new_n1832;
  assign new_n2269 = ~new_n2267 & ~new_n2268;
  assign new_n2270 = new_n1842 & ~new_n2269;
  assign new_n2271 = ~new_n2266 & ~new_n2270;
  assign new_n2272 = new_n1855 & ~new_n2271;
  assign new_n2273 = ~new_n2265 & ~new_n2272;
  assign new_n2274 = new_n1869 & ~new_n2273;
  assign new_n2275 = ~new_n1756 & new_n2274;
  assign new_n2276 = new_n364 & new_n2275;
  assign new_n2277 = ~new_n364 & ~new_n2275;
  assign new_n2278 = ~new_n2276 & ~new_n2277;
  assign new_n2279 = ~new_n2264 & ~new_n2278;
  assign new_n2280 = new_n2250 & new_n2279;
  assign new_n2281 = ~new_n2221 & new_n2280;
  assign new_n2282 = ~new_n383 & new_n2232;
  assign new_n2283 = ~new_n2249 & new_n2282;
  assign new_n2284 = ~new_n377 & new_n2246;
  assign new_n2285 = ~new_n2283 & ~new_n2284;
  assign new_n2286 = new_n2279 & ~new_n2285;
  assign new_n2287 = ~new_n370 & new_n2261;
  assign new_n2288 = ~new_n2278 & new_n2287;
  assign new_n2289 = ~new_n364 & new_n2275;
  assign new_n2290 = ~new_n2288 & ~new_n2289;
  assign new_n2291 = ~new_n2286 & new_n2290;
  assign new_n2292 = ~new_n2281 & new_n2291;
  assign new_n2293 = ~new_n1869 & new_n2174;
  assign new_n2294 = ~new_n1855 & ~new_n2228;
  assign new_n2295 = ~new_n1842 & ~new_n2255;
  assign new_n2296 = ~new_n1765 & ~new_n1832;
  assign new_n2297 = new_n1842 & new_n2296;
  assign new_n2298 = ~new_n2295 & ~new_n2297;
  assign new_n2299 = new_n1855 & ~new_n2298;
  assign new_n2300 = ~new_n2294 & ~new_n2299;
  assign new_n2301 = new_n1869 & ~new_n2300;
  assign new_n2302 = ~new_n2293 & ~new_n2301;
  assign new_n2303 = ~new_n1756 & ~new_n2302;
  assign new_n2304 = new_n355 & new_n2303;
  assign new_n2305 = ~new_n355 & ~new_n2303;
  assign new_n2306 = ~new_n2304 & ~new_n2305;
  assign new_n2307 = ~new_n1869 & new_n2182;
  assign new_n2308 = ~new_n1855 & ~new_n2242;
  assign new_n2309 = ~new_n1842 & ~new_n2269;
  assign new_n2310 = new_n1855 & new_n2309;
  assign new_n2311 = ~new_n2308 & ~new_n2310;
  assign new_n2312 = new_n1869 & ~new_n2311;
  assign new_n2313 = ~new_n2307 & ~new_n2312;
  assign new_n2314 = ~new_n1756 & ~new_n2313;
  assign new_n2315 = new_n349 & new_n2314;
  assign new_n2316 = ~new_n349 & ~new_n2314;
  assign new_n2317 = ~new_n2315 & ~new_n2316;
  assign new_n2318 = ~new_n2306 & ~new_n2317;
  assign new_n2319 = ~new_n1869 & new_n2197;
  assign new_n2320 = ~new_n1855 & ~new_n2257;
  assign new_n2321 = ~new_n1842 & new_n2296;
  assign new_n2322 = new_n1855 & new_n2321;
  assign new_n2323 = ~new_n2320 & ~new_n2322;
  assign new_n2324 = new_n1869 & ~new_n2323;
  assign new_n2325 = ~new_n2319 & ~new_n2324;
  assign new_n2326 = ~new_n1756 & ~new_n2325;
  assign new_n2327 = new_n342 & new_n2326;
  assign new_n2328 = ~new_n342 & ~new_n2326;
  assign new_n2329 = ~new_n2327 & ~new_n2328;
  assign new_n2330 = ~new_n1869 & new_n2209;
  assign new_n2331 = ~new_n1855 & ~new_n2271;
  assign new_n2332 = new_n1869 & new_n2331;
  assign new_n2333 = ~new_n2330 & ~new_n2332;
  assign new_n2334 = ~new_n1756 & ~new_n2333;
  assign new_n2335 = new_n336 & new_n2334;
  assign new_n2336 = ~new_n336 & ~new_n2334;
  assign new_n2337 = ~new_n2335 & ~new_n2336;
  assign new_n2338 = ~new_n2329 & ~new_n2337;
  assign new_n2339 = new_n2318 & new_n2338;
  assign new_n2340 = ~new_n2292 & new_n2339;
  assign new_n2341 = ~new_n355 & new_n2303;
  assign new_n2342 = ~new_n2317 & new_n2341;
  assign new_n2343 = ~new_n349 & new_n2314;
  assign new_n2344 = ~new_n2342 & ~new_n2343;
  assign new_n2345 = new_n2338 & ~new_n2344;
  assign new_n2346 = ~new_n342 & new_n2326;
  assign new_n2347 = ~new_n2337 & new_n2346;
  assign new_n2348 = ~new_n336 & new_n2334;
  assign new_n2349 = ~new_n2347 & ~new_n2348;
  assign new_n2350 = ~new_n2345 & new_n2349;
  assign new_n2351 = ~new_n2340 & new_n2350;
  assign new_n2352 = ~new_n1869 & ~new_n2230;
  assign new_n2353 = ~new_n1855 & ~new_n2298;
  assign new_n2354 = new_n1869 & new_n2353;
  assign new_n2355 = ~new_n2352 & ~new_n2354;
  assign new_n2356 = ~new_n1756 & ~new_n2355;
  assign new_n2357 = new_n328 & new_n2356;
  assign new_n2358 = ~new_n328 & ~new_n2356;
  assign new_n2359 = ~new_n2357 & ~new_n2358;
  assign new_n2360 = ~new_n1869 & ~new_n2244;
  assign new_n2361 = ~new_n1855 & new_n2309;
  assign new_n2362 = new_n1869 & new_n2361;
  assign new_n2363 = ~new_n2360 & ~new_n2362;
  assign new_n2364 = ~new_n1756 & ~new_n2363;
  assign new_n2365 = new_n322 & new_n2364;
  assign new_n2366 = ~new_n322 & ~new_n2364;
  assign new_n2367 = ~new_n2365 & ~new_n2366;
  assign new_n2368 = ~new_n2359 & ~new_n2367;
  assign new_n2369 = ~new_n2351 & new_n2368;
  assign new_n2370 = ~new_n328 & new_n2356;
  assign new_n2371 = ~new_n2367 & new_n2370;
  assign new_n2372 = ~new_n322 & new_n2364;
  assign new_n2373 = ~new_n2371 & ~new_n2372;
  assign new_n2374 = ~new_n2369 & new_n2373;
  assign new_n2375 = ~new_n1869 & ~new_n2259;
  assign new_n2376 = ~new_n1855 & new_n2321;
  assign new_n2377 = new_n1869 & new_n2376;
  assign new_n2378 = ~new_n2375 & ~new_n2377;
  assign new_n2379 = ~new_n1756 & ~new_n2378;
  assign new_n2380 = new_n315 & new_n2379;
  assign new_n2381 = ~new_n315 & ~new_n2379;
  assign new_n2382 = ~new_n2380 & ~new_n2381;
  assign new_n2383 = ~new_n2374 & ~new_n2382;
  assign new_n2384 = ~new_n315 & new_n2379;
  assign new_n2385 = ~new_n2383 & ~new_n2384;
  assign new_n2386 = ~new_n1869 & ~new_n2273;
  assign new_n2387 = ~new_n1756 & new_n2386;
  assign new_n2388 = new_n309 & new_n2387;
  assign new_n2389 = ~new_n309 & ~new_n2387;
  assign new_n2390 = ~new_n2388 & ~new_n2389;
  assign new_n2391 = new_n2385 & ~new_n2390;
  assign new_n2392 = ~new_n2385 & new_n2390;
  assign new_n2393 = ~new_n2391 & ~new_n2392;
  assign new_n2394 = ~new_n1794 & ~new_n2393;
  assign new_n2395 = new_n1727 & new_n2394;
  assign new_n2396 = ~new_n2171 & ~new_n2395;
  assign new_n2397 = lo33 & ~new_n1700;
  assign new_n2398 = ~lo02 & lo76;
  assign new_n2399 = ~lo03 & new_n2398;
  assign new_n2400 = ~lo04 & new_n2399;
  assign new_n2401 = ~lo05 & new_n2400;
  assign new_n2402 = lo35 & new_n2401;
  assign new_n2403 = lo18 & new_n2402;
  assign new_n2404 = lo02 & lo76;
  assign new_n2405 = ~lo02 & lo77;
  assign new_n2406 = ~new_n2404 & ~new_n2405;
  assign new_n2407 = ~lo03 & ~new_n2406;
  assign new_n2408 = ~lo04 & new_n2407;
  assign new_n2409 = ~lo05 & new_n2408;
  assign new_n2410 = lo35 & new_n2409;
  assign new_n2411 = ~lo19 & new_n2410;
  assign new_n2412 = lo19 & ~new_n2410;
  assign new_n2413 = ~new_n2411 & ~new_n2412;
  assign new_n2414 = new_n2403 & ~new_n2413;
  assign new_n2415 = lo19 & new_n2410;
  assign new_n2416 = ~new_n2414 & ~new_n2415;
  assign new_n2417 = lo03 & new_n2398;
  assign new_n2418 = lo02 & lo77;
  assign new_n2419 = ~lo02 & lo78;
  assign new_n2420 = ~new_n2418 & ~new_n2419;
  assign new_n2421 = ~lo03 & ~new_n2420;
  assign new_n2422 = ~new_n2417 & ~new_n2421;
  assign new_n2423 = ~lo04 & ~new_n2422;
  assign new_n2424 = ~lo05 & new_n2423;
  assign new_n2425 = lo35 & new_n2424;
  assign new_n2426 = ~lo20 & new_n2425;
  assign new_n2427 = lo20 & ~new_n2425;
  assign new_n2428 = ~new_n2426 & ~new_n2427;
  assign new_n2429 = lo03 & ~new_n2406;
  assign new_n2430 = lo02 & lo78;
  assign new_n2431 = ~lo02 & lo79;
  assign new_n2432 = ~new_n2430 & ~new_n2431;
  assign new_n2433 = ~lo03 & ~new_n2432;
  assign new_n2434 = ~new_n2429 & ~new_n2433;
  assign new_n2435 = ~lo04 & ~new_n2434;
  assign new_n2436 = ~lo05 & new_n2435;
  assign new_n2437 = lo35 & new_n2436;
  assign new_n2438 = ~lo21 & new_n2437;
  assign new_n2439 = lo21 & ~new_n2437;
  assign new_n2440 = ~new_n2438 & ~new_n2439;
  assign new_n2441 = ~new_n2428 & ~new_n2440;
  assign new_n2442 = ~new_n2416 & new_n2441;
  assign new_n2443 = lo20 & new_n2425;
  assign new_n2444 = ~new_n2440 & new_n2443;
  assign new_n2445 = lo21 & new_n2437;
  assign new_n2446 = ~new_n2444 & ~new_n2445;
  assign new_n2447 = ~new_n2442 & new_n2446;
  assign new_n2448 = lo04 & new_n2399;
  assign new_n2449 = lo03 & ~new_n2420;
  assign new_n2450 = lo02 & lo79;
  assign new_n2451 = ~lo02 & lo80;
  assign new_n2452 = ~new_n2450 & ~new_n2451;
  assign new_n2453 = ~lo03 & ~new_n2452;
  assign new_n2454 = ~new_n2449 & ~new_n2453;
  assign new_n2455 = ~lo04 & ~new_n2454;
  assign new_n2456 = ~new_n2448 & ~new_n2455;
  assign new_n2457 = ~lo05 & ~new_n2456;
  assign new_n2458 = lo35 & new_n2457;
  assign new_n2459 = ~lo22 & new_n2458;
  assign new_n2460 = lo22 & ~new_n2458;
  assign new_n2461 = ~new_n2459 & ~new_n2460;
  assign new_n2462 = lo04 & new_n2407;
  assign new_n2463 = lo03 & ~new_n2432;
  assign new_n2464 = lo02 & lo80;
  assign new_n2465 = ~lo02 & lo81;
  assign new_n2466 = ~new_n2464 & ~new_n2465;
  assign new_n2467 = ~lo03 & ~new_n2466;
  assign new_n2468 = ~new_n2463 & ~new_n2467;
  assign new_n2469 = ~lo04 & ~new_n2468;
  assign new_n2470 = ~new_n2462 & ~new_n2469;
  assign new_n2471 = ~lo05 & ~new_n2470;
  assign new_n2472 = lo35 & new_n2471;
  assign new_n2473 = ~lo23 & new_n2472;
  assign new_n2474 = lo23 & ~new_n2472;
  assign new_n2475 = ~new_n2473 & ~new_n2474;
  assign new_n2476 = ~new_n2461 & ~new_n2475;
  assign new_n2477 = lo04 & ~new_n2422;
  assign new_n2478 = lo03 & ~new_n2452;
  assign new_n2479 = lo02 & lo81;
  assign new_n2480 = ~lo02 & lo82;
  assign new_n2481 = ~new_n2479 & ~new_n2480;
  assign new_n2482 = ~lo03 & ~new_n2481;
  assign new_n2483 = ~new_n2478 & ~new_n2482;
  assign new_n2484 = ~lo04 & ~new_n2483;
  assign new_n2485 = ~new_n2477 & ~new_n2484;
  assign new_n2486 = ~lo05 & ~new_n2485;
  assign new_n2487 = lo35 & new_n2486;
  assign new_n2488 = ~lo24 & new_n2487;
  assign new_n2489 = lo24 & ~new_n2487;
  assign new_n2490 = ~new_n2488 & ~new_n2489;
  assign new_n2491 = lo04 & ~new_n2434;
  assign new_n2492 = lo03 & ~new_n2466;
  assign new_n2493 = lo02 & lo82;
  assign new_n2494 = ~lo02 & lo83;
  assign new_n2495 = ~new_n2493 & ~new_n2494;
  assign new_n2496 = ~lo03 & ~new_n2495;
  assign new_n2497 = ~new_n2492 & ~new_n2496;
  assign new_n2498 = ~lo04 & ~new_n2497;
  assign new_n2499 = ~new_n2491 & ~new_n2498;
  assign new_n2500 = ~lo05 & ~new_n2499;
  assign new_n2501 = lo35 & new_n2500;
  assign new_n2502 = ~lo25 & new_n2501;
  assign new_n2503 = lo25 & ~new_n2501;
  assign new_n2504 = ~new_n2502 & ~new_n2503;
  assign new_n2505 = ~new_n2490 & ~new_n2504;
  assign new_n2506 = new_n2476 & new_n2505;
  assign new_n2507 = ~new_n2447 & new_n2506;
  assign new_n2508 = lo22 & new_n2458;
  assign new_n2509 = ~new_n2475 & new_n2508;
  assign new_n2510 = lo23 & new_n2472;
  assign new_n2511 = ~new_n2509 & ~new_n2510;
  assign new_n2512 = new_n2505 & ~new_n2511;
  assign new_n2513 = lo24 & new_n2487;
  assign new_n2514 = ~new_n2504 & new_n2513;
  assign new_n2515 = lo25 & new_n2501;
  assign new_n2516 = ~new_n2514 & ~new_n2515;
  assign new_n2517 = ~new_n2512 & new_n2516;
  assign new_n2518 = ~new_n2507 & new_n2517;
  assign new_n2519 = lo05 & new_n2400;
  assign new_n2520 = lo04 & ~new_n2454;
  assign new_n2521 = lo03 & ~new_n2481;
  assign new_n2522 = lo02 & lo83;
  assign new_n2523 = ~lo03 & new_n2522;
  assign new_n2524 = ~new_n2521 & ~new_n2523;
  assign new_n2525 = ~lo04 & ~new_n2524;
  assign new_n2526 = ~new_n2520 & ~new_n2525;
  assign new_n2527 = ~lo05 & ~new_n2526;
  assign new_n2528 = ~new_n2519 & ~new_n2527;
  assign new_n2529 = lo35 & ~new_n2528;
  assign new_n2530 = ~lo26 & new_n2529;
  assign new_n2531 = lo26 & ~new_n2529;
  assign new_n2532 = ~new_n2530 & ~new_n2531;
  assign new_n2533 = lo05 & new_n2408;
  assign new_n2534 = lo04 & ~new_n2468;
  assign new_n2535 = lo03 & ~new_n2495;
  assign new_n2536 = ~lo04 & new_n2535;
  assign new_n2537 = ~new_n2534 & ~new_n2536;
  assign new_n2538 = ~lo05 & ~new_n2537;
  assign new_n2539 = ~new_n2533 & ~new_n2538;
  assign new_n2540 = lo35 & ~new_n2539;
  assign new_n2541 = ~lo27 & new_n2540;
  assign new_n2542 = lo27 & ~new_n2540;
  assign new_n2543 = ~new_n2541 & ~new_n2542;
  assign new_n2544 = ~new_n2532 & ~new_n2543;
  assign new_n2545 = lo05 & new_n2423;
  assign new_n2546 = lo04 & ~new_n2483;
  assign new_n2547 = lo03 & new_n2522;
  assign new_n2548 = ~lo04 & new_n2547;
  assign new_n2549 = ~new_n2546 & ~new_n2548;
  assign new_n2550 = ~lo05 & ~new_n2549;
  assign new_n2551 = ~new_n2545 & ~new_n2550;
  assign new_n2552 = lo35 & ~new_n2551;
  assign new_n2553 = ~lo28 & new_n2552;
  assign new_n2554 = lo28 & ~new_n2552;
  assign new_n2555 = ~new_n2553 & ~new_n2554;
  assign new_n2556 = lo05 & new_n2435;
  assign new_n2557 = lo04 & ~new_n2497;
  assign new_n2558 = ~lo05 & new_n2557;
  assign new_n2559 = ~new_n2556 & ~new_n2558;
  assign new_n2560 = lo35 & ~new_n2559;
  assign new_n2561 = ~lo29 & new_n2560;
  assign new_n2562 = lo29 & ~new_n2560;
  assign new_n2563 = ~new_n2561 & ~new_n2562;
  assign new_n2564 = ~new_n2555 & ~new_n2563;
  assign new_n2565 = new_n2544 & new_n2564;
  assign new_n2566 = ~new_n2518 & new_n2565;
  assign new_n2567 = lo26 & new_n2529;
  assign new_n2568 = ~new_n2543 & new_n2567;
  assign new_n2569 = lo27 & new_n2540;
  assign new_n2570 = ~new_n2568 & ~new_n2569;
  assign new_n2571 = new_n2564 & ~new_n2570;
  assign new_n2572 = lo28 & new_n2552;
  assign new_n2573 = ~new_n2563 & new_n2572;
  assign new_n2574 = lo29 & new_n2560;
  assign new_n2575 = ~new_n2573 & ~new_n2574;
  assign new_n2576 = ~new_n2571 & new_n2575;
  assign new_n2577 = ~new_n2566 & new_n2576;
  assign new_n2578 = lo05 & ~new_n2456;
  assign new_n2579 = lo04 & ~new_n2524;
  assign new_n2580 = ~lo05 & new_n2579;
  assign new_n2581 = ~new_n2578 & ~new_n2580;
  assign new_n2582 = lo35 & ~new_n2581;
  assign new_n2583 = ~lo30 & new_n2582;
  assign new_n2584 = lo30 & ~new_n2582;
  assign new_n2585 = ~new_n2583 & ~new_n2584;
  assign new_n2586 = lo05 & ~new_n2470;
  assign new_n2587 = lo04 & new_n2535;
  assign new_n2588 = ~lo05 & new_n2587;
  assign new_n2589 = ~new_n2586 & ~new_n2588;
  assign new_n2590 = lo35 & ~new_n2589;
  assign new_n2591 = ~lo31 & new_n2590;
  assign new_n2592 = lo31 & ~new_n2590;
  assign new_n2593 = ~new_n2591 & ~new_n2592;
  assign new_n2594 = ~new_n2585 & ~new_n2593;
  assign new_n2595 = ~new_n2577 & new_n2594;
  assign new_n2596 = lo30 & new_n2582;
  assign new_n2597 = ~new_n2593 & new_n2596;
  assign new_n2598 = lo31 & new_n2590;
  assign new_n2599 = ~new_n2597 & ~new_n2598;
  assign new_n2600 = ~new_n2595 & new_n2599;
  assign new_n2601 = lo05 & ~new_n2485;
  assign new_n2602 = lo04 & new_n2547;
  assign new_n2603 = ~lo05 & new_n2602;
  assign new_n2604 = ~new_n2601 & ~new_n2603;
  assign new_n2605 = lo35 & ~new_n2604;
  assign new_n2606 = ~lo32 & new_n2605;
  assign new_n2607 = lo32 & ~new_n2605;
  assign new_n2608 = ~new_n2606 & ~new_n2607;
  assign new_n2609 = ~new_n2600 & ~new_n2608;
  assign new_n2610 = lo32 & new_n2605;
  assign new_n2611 = ~new_n2609 & ~new_n2610;
  assign new_n2612 = lo05 & ~new_n2499;
  assign new_n2613 = lo35 & new_n2612;
  assign new_n2614 = ~lo33 & new_n2613;
  assign new_n2615 = lo33 & ~new_n2613;
  assign new_n2616 = ~new_n2614 & ~new_n2615;
  assign new_n2617 = new_n2611 & ~new_n2616;
  assign new_n2618 = ~new_n2611 & new_n2616;
  assign new_n2619 = ~new_n2617 & ~new_n2618;
  assign new_n2620 = lo43 & ~new_n2619;
  assign new_n2621 = new_n1700 & new_n2620;
  assign li33 = new_n2397 | new_n2621;
  assign new_n2623 = new_n2396 & li33;
  assign new_n2624 = ~new_n2396 & ~li33;
  assign new_n2625 = ~new_n2623 & ~new_n2624;
  assign new_n2626 = ~new_n315 & ~new_n1727;
  assign new_n2627 = new_n2374 & ~new_n2382;
  assign new_n2628 = ~new_n2374 & new_n2382;
  assign new_n2629 = ~new_n2627 & ~new_n2628;
  assign new_n2630 = ~new_n1794 & ~new_n2629;
  assign new_n2631 = new_n1727 & new_n2630;
  assign new_n2632 = ~new_n2626 & ~new_n2631;
  assign new_n2633 = lo32 & ~new_n1700;
  assign new_n2634 = new_n2600 & ~new_n2608;
  assign new_n2635 = ~new_n2600 & new_n2608;
  assign new_n2636 = ~new_n2634 & ~new_n2635;
  assign new_n2637 = lo43 & ~new_n2636;
  assign new_n2638 = new_n1700 & new_n2637;
  assign li32 = new_n2633 | new_n2638;
  assign new_n2640 = new_n2632 & li32;
  assign new_n2641 = ~new_n2632 & ~li32;
  assign new_n2642 = ~new_n2640 & ~new_n2641;
  assign new_n2643 = new_n2625 & new_n2642;
  assign new_n2644 = ~new_n322 & ~new_n1727;
  assign new_n2645 = ~new_n2351 & ~new_n2359;
  assign new_n2646 = ~new_n2370 & ~new_n2645;
  assign new_n2647 = ~new_n2367 & new_n2646;
  assign new_n2648 = new_n2367 & ~new_n2646;
  assign new_n2649 = ~new_n2647 & ~new_n2648;
  assign new_n2650 = ~new_n1794 & ~new_n2649;
  assign new_n2651 = new_n1727 & new_n2650;
  assign new_n2652 = ~new_n2644 & ~new_n2651;
  assign new_n2653 = lo31 & ~new_n1700;
  assign new_n2654 = ~new_n2577 & ~new_n2585;
  assign new_n2655 = ~new_n2596 & ~new_n2654;
  assign new_n2656 = ~new_n2593 & new_n2655;
  assign new_n2657 = new_n2593 & ~new_n2655;
  assign new_n2658 = ~new_n2656 & ~new_n2657;
  assign new_n2659 = lo43 & ~new_n2658;
  assign new_n2660 = new_n1700 & new_n2659;
  assign li31 = new_n2653 | new_n2660;
  assign new_n2662 = new_n2652 & li31;
  assign new_n2663 = ~new_n2652 & ~li31;
  assign new_n2664 = ~new_n2662 & ~new_n2663;
  assign new_n2665 = ~new_n328 & ~new_n1727;
  assign new_n2666 = new_n2351 & ~new_n2359;
  assign new_n2667 = ~new_n2351 & new_n2359;
  assign new_n2668 = ~new_n2666 & ~new_n2667;
  assign new_n2669 = ~new_n1794 & ~new_n2668;
  assign new_n2670 = new_n1727 & new_n2669;
  assign new_n2671 = ~new_n2665 & ~new_n2670;
  assign new_n2672 = lo30 & ~new_n1700;
  assign new_n2673 = new_n2577 & ~new_n2585;
  assign new_n2674 = ~new_n2577 & new_n2585;
  assign new_n2675 = ~new_n2673 & ~new_n2674;
  assign new_n2676 = lo43 & ~new_n2675;
  assign new_n2677 = new_n1700 & new_n2676;
  assign li30 = new_n2672 | new_n2677;
  assign new_n2679 = new_n2671 & li30;
  assign new_n2680 = ~new_n2671 & ~li30;
  assign new_n2681 = ~new_n2679 & ~new_n2680;
  assign new_n2682 = new_n2664 & new_n2681;
  assign new_n2683 = new_n2643 & new_n2682;
  assign new_n2684 = ~new_n336 & ~new_n1727;
  assign new_n2685 = ~new_n2292 & new_n2318;
  assign new_n2686 = new_n2344 & ~new_n2685;
  assign new_n2687 = ~new_n2329 & ~new_n2686;
  assign new_n2688 = ~new_n2346 & ~new_n2687;
  assign new_n2689 = ~new_n2337 & new_n2688;
  assign new_n2690 = new_n2337 & ~new_n2688;
  assign new_n2691 = ~new_n2689 & ~new_n2690;
  assign new_n2692 = ~new_n1794 & ~new_n2691;
  assign new_n2693 = new_n1727 & new_n2692;
  assign new_n2694 = ~new_n2684 & ~new_n2693;
  assign new_n2695 = lo29 & ~new_n1700;
  assign new_n2696 = ~new_n2518 & new_n2544;
  assign new_n2697 = new_n2570 & ~new_n2696;
  assign new_n2698 = ~new_n2555 & ~new_n2697;
  assign new_n2699 = ~new_n2572 & ~new_n2698;
  assign new_n2700 = ~new_n2563 & new_n2699;
  assign new_n2701 = new_n2563 & ~new_n2699;
  assign new_n2702 = ~new_n2700 & ~new_n2701;
  assign new_n2703 = lo43 & ~new_n2702;
  assign new_n2704 = new_n1700 & new_n2703;
  assign li29 = new_n2695 | new_n2704;
  assign new_n2706 = new_n2694 & li29;
  assign new_n2707 = ~new_n2694 & ~li29;
  assign new_n2708 = ~new_n2706 & ~new_n2707;
  assign new_n2709 = ~new_n342 & ~new_n1727;
  assign new_n2710 = ~new_n2329 & new_n2686;
  assign new_n2711 = new_n2329 & ~new_n2686;
  assign new_n2712 = ~new_n2710 & ~new_n2711;
  assign new_n2713 = ~new_n1794 & ~new_n2712;
  assign new_n2714 = new_n1727 & new_n2713;
  assign new_n2715 = ~new_n2709 & ~new_n2714;
  assign new_n2716 = lo28 & ~new_n1700;
  assign new_n2717 = ~new_n2555 & new_n2697;
  assign new_n2718 = new_n2555 & ~new_n2697;
  assign new_n2719 = ~new_n2717 & ~new_n2718;
  assign new_n2720 = lo43 & ~new_n2719;
  assign new_n2721 = new_n1700 & new_n2720;
  assign li28 = new_n2716 | new_n2721;
  assign new_n2723 = new_n2715 & li28;
  assign new_n2724 = ~new_n2715 & ~li28;
  assign new_n2725 = ~new_n2723 & ~new_n2724;
  assign new_n2726 = new_n2708 & new_n2725;
  assign new_n2727 = ~new_n349 & ~new_n1727;
  assign new_n2728 = ~new_n2292 & ~new_n2306;
  assign new_n2729 = ~new_n2341 & ~new_n2728;
  assign new_n2730 = ~new_n2317 & new_n2729;
  assign new_n2731 = new_n2317 & ~new_n2729;
  assign new_n2732 = ~new_n2730 & ~new_n2731;
  assign new_n2733 = ~new_n1794 & ~new_n2732;
  assign new_n2734 = new_n1727 & new_n2733;
  assign new_n2735 = ~new_n2727 & ~new_n2734;
  assign new_n2736 = lo27 & ~new_n1700;
  assign new_n2737 = ~new_n2518 & ~new_n2532;
  assign new_n2738 = ~new_n2567 & ~new_n2737;
  assign new_n2739 = ~new_n2543 & new_n2738;
  assign new_n2740 = new_n2543 & ~new_n2738;
  assign new_n2741 = ~new_n2739 & ~new_n2740;
  assign new_n2742 = lo43 & ~new_n2741;
  assign new_n2743 = new_n1700 & new_n2742;
  assign li27 = new_n2736 | new_n2743;
  assign new_n2745 = new_n2735 & li27;
  assign new_n2746 = ~new_n2735 & ~li27;
  assign new_n2747 = ~new_n2745 & ~new_n2746;
  assign new_n2748 = ~new_n355 & ~new_n1727;
  assign new_n2749 = new_n2292 & ~new_n2306;
  assign new_n2750 = ~new_n2292 & new_n2306;
  assign new_n2751 = ~new_n2749 & ~new_n2750;
  assign new_n2752 = ~new_n1794 & ~new_n2751;
  assign new_n2753 = new_n1727 & new_n2752;
  assign new_n2754 = ~new_n2748 & ~new_n2753;
  assign new_n2755 = lo26 & ~new_n1700;
  assign new_n2756 = new_n2518 & ~new_n2532;
  assign new_n2757 = ~new_n2518 & new_n2532;
  assign new_n2758 = ~new_n2756 & ~new_n2757;
  assign new_n2759 = lo43 & ~new_n2758;
  assign new_n2760 = new_n1700 & new_n2759;
  assign li26 = new_n2755 | new_n2760;
  assign new_n2762 = new_n2754 & li26;
  assign new_n2763 = ~new_n2754 & ~li26;
  assign new_n2764 = ~new_n2762 & ~new_n2763;
  assign new_n2765 = new_n2747 & new_n2764;
  assign new_n2766 = new_n2726 & new_n2765;
  assign new_n2767 = new_n2683 & new_n2766;
  assign new_n2768 = ~new_n364 & ~new_n1727;
  assign new_n2769 = ~new_n2221 & new_n2250;
  assign new_n2770 = new_n2285 & ~new_n2769;
  assign new_n2771 = ~new_n2264 & ~new_n2770;
  assign new_n2772 = ~new_n2287 & ~new_n2771;
  assign new_n2773 = ~new_n2278 & new_n2772;
  assign new_n2774 = new_n2278 & ~new_n2772;
  assign new_n2775 = ~new_n2773 & ~new_n2774;
  assign new_n2776 = ~new_n1794 & ~new_n2775;
  assign new_n2777 = new_n1727 & new_n2776;
  assign new_n2778 = ~new_n2768 & ~new_n2777;
  assign new_n2779 = lo25 & ~new_n1700;
  assign new_n2780 = ~new_n2447 & new_n2476;
  assign new_n2781 = new_n2511 & ~new_n2780;
  assign new_n2782 = ~new_n2490 & ~new_n2781;
  assign new_n2783 = ~new_n2513 & ~new_n2782;
  assign new_n2784 = ~new_n2504 & new_n2783;
  assign new_n2785 = new_n2504 & ~new_n2783;
  assign new_n2786 = ~new_n2784 & ~new_n2785;
  assign new_n2787 = lo43 & ~new_n2786;
  assign new_n2788 = new_n1700 & new_n2787;
  assign li25 = new_n2779 | new_n2788;
  assign new_n2790 = new_n2778 & li25;
  assign new_n2791 = ~new_n2778 & ~li25;
  assign new_n2792 = ~new_n2790 & ~new_n2791;
  assign new_n2793 = ~new_n370 & ~new_n1727;
  assign new_n2794 = ~new_n2264 & new_n2770;
  assign new_n2795 = new_n2264 & ~new_n2770;
  assign new_n2796 = ~new_n2794 & ~new_n2795;
  assign new_n2797 = ~new_n1794 & ~new_n2796;
  assign new_n2798 = new_n1727 & new_n2797;
  assign new_n2799 = ~new_n2793 & ~new_n2798;
  assign new_n2800 = lo24 & ~new_n1700;
  assign new_n2801 = ~new_n2490 & new_n2781;
  assign new_n2802 = new_n2490 & ~new_n2781;
  assign new_n2803 = ~new_n2801 & ~new_n2802;
  assign new_n2804 = lo43 & ~new_n2803;
  assign new_n2805 = new_n1700 & new_n2804;
  assign li24 = new_n2800 | new_n2805;
  assign new_n2807 = new_n2799 & li24;
  assign new_n2808 = ~new_n2799 & ~li24;
  assign new_n2809 = ~new_n2807 & ~new_n2808;
  assign new_n2810 = new_n2792 & new_n2809;
  assign new_n2811 = ~new_n377 & ~new_n1727;
  assign new_n2812 = ~new_n2221 & ~new_n2235;
  assign new_n2813 = ~new_n2282 & ~new_n2812;
  assign new_n2814 = ~new_n2249 & new_n2813;
  assign new_n2815 = new_n2249 & ~new_n2813;
  assign new_n2816 = ~new_n2814 & ~new_n2815;
  assign new_n2817 = ~new_n1794 & ~new_n2816;
  assign new_n2818 = new_n1727 & new_n2817;
  assign new_n2819 = ~new_n2811 & ~new_n2818;
  assign new_n2820 = lo23 & ~new_n1700;
  assign new_n2821 = ~new_n2447 & ~new_n2461;
  assign new_n2822 = ~new_n2508 & ~new_n2821;
  assign new_n2823 = ~new_n2475 & new_n2822;
  assign new_n2824 = new_n2475 & ~new_n2822;
  assign new_n2825 = ~new_n2823 & ~new_n2824;
  assign new_n2826 = lo43 & ~new_n2825;
  assign new_n2827 = new_n1700 & new_n2826;
  assign li23 = new_n2820 | new_n2827;
  assign new_n2829 = new_n2819 & li23;
  assign new_n2830 = ~new_n2819 & ~li23;
  assign new_n2831 = ~new_n2829 & ~new_n2830;
  assign new_n2832 = ~new_n383 & ~new_n1727;
  assign new_n2833 = new_n2221 & ~new_n2235;
  assign new_n2834 = ~new_n2221 & new_n2235;
  assign new_n2835 = ~new_n2833 & ~new_n2834;
  assign new_n2836 = ~new_n1794 & ~new_n2835;
  assign new_n2837 = new_n1727 & new_n2836;
  assign new_n2838 = ~new_n2832 & ~new_n2837;
  assign new_n2839 = lo22 & ~new_n1700;
  assign new_n2840 = new_n2447 & ~new_n2461;
  assign new_n2841 = ~new_n2447 & new_n2461;
  assign new_n2842 = ~new_n2840 & ~new_n2841;
  assign new_n2843 = lo43 & ~new_n2842;
  assign new_n2844 = new_n1700 & new_n2843;
  assign li22 = new_n2839 | new_n2844;
  assign new_n2846 = new_n2838 & li22;
  assign new_n2847 = ~new_n2838 & ~li22;
  assign new_n2848 = ~new_n2846 & ~new_n2847;
  assign new_n2849 = new_n2831 & new_n2848;
  assign new_n2850 = new_n2810 & new_n2849;
  assign new_n2851 = ~new_n391 & ~new_n1727;
  assign new_n2852 = ~new_n2190 & ~new_n2202;
  assign new_n2853 = ~new_n2217 & ~new_n2852;
  assign new_n2854 = ~new_n2214 & new_n2853;
  assign new_n2855 = new_n2214 & ~new_n2853;
  assign new_n2856 = ~new_n2854 & ~new_n2855;
  assign new_n2857 = ~new_n1794 & ~new_n2856;
  assign new_n2858 = new_n1727 & new_n2857;
  assign new_n2859 = ~new_n2851 & ~new_n2858;
  assign new_n2860 = lo21 & ~new_n1700;
  assign new_n2861 = ~new_n2416 & ~new_n2428;
  assign new_n2862 = ~new_n2443 & ~new_n2861;
  assign new_n2863 = ~new_n2440 & new_n2862;
  assign new_n2864 = new_n2440 & ~new_n2862;
  assign new_n2865 = ~new_n2863 & ~new_n2864;
  assign new_n2866 = lo43 & ~new_n2865;
  assign new_n2867 = new_n1700 & new_n2866;
  assign li21 = new_n2860 | new_n2867;
  assign new_n2869 = new_n2859 & li21;
  assign new_n2870 = ~new_n2859 & ~li21;
  assign new_n2871 = ~new_n2869 & ~new_n2870;
  assign new_n2872 = ~new_n397 & ~new_n1727;
  assign new_n2873 = new_n2190 & ~new_n2202;
  assign new_n2874 = ~new_n2190 & new_n2202;
  assign new_n2875 = ~new_n2873 & ~new_n2874;
  assign new_n2876 = ~new_n1794 & ~new_n2875;
  assign new_n2877 = new_n1727 & new_n2876;
  assign new_n2878 = ~new_n2872 & ~new_n2877;
  assign new_n2879 = lo20 & ~new_n1700;
  assign new_n2880 = new_n2416 & ~new_n2428;
  assign new_n2881 = ~new_n2416 & new_n2428;
  assign new_n2882 = ~new_n2880 & ~new_n2881;
  assign new_n2883 = lo43 & ~new_n2882;
  assign new_n2884 = new_n1700 & new_n2883;
  assign li20 = new_n2879 | new_n2884;
  assign new_n2886 = new_n2878 & li20;
  assign new_n2887 = ~new_n2878 & ~li20;
  assign new_n2888 = ~new_n2886 & ~new_n2887;
  assign new_n2889 = new_n2871 & new_n2888;
  assign new_n2890 = ~new_n404 & ~new_n1727;
  assign new_n2891 = ~new_n2177 & ~new_n2187;
  assign new_n2892 = new_n2177 & new_n2187;
  assign new_n2893 = ~new_n2891 & ~new_n2892;
  assign new_n2894 = ~new_n1794 & ~new_n2893;
  assign new_n2895 = new_n1727 & new_n2894;
  assign new_n2896 = ~new_n2890 & ~new_n2895;
  assign new_n2897 = lo19 & ~new_n1700;
  assign new_n2898 = ~new_n2403 & ~new_n2413;
  assign new_n2899 = new_n2403 & new_n2413;
  assign new_n2900 = ~new_n2898 & ~new_n2899;
  assign new_n2901 = lo43 & ~new_n2900;
  assign new_n2902 = new_n1700 & new_n2901;
  assign li19 = new_n2897 | new_n2902;
  assign new_n2904 = new_n2896 & li19;
  assign new_n2905 = ~new_n2896 & ~li19;
  assign new_n2906 = ~new_n2904 & ~new_n2905;
  assign new_n2907 = ~new_n410 & ~new_n1727;
  assign new_n2908 = new_n410 & new_n2176;
  assign new_n2909 = ~new_n410 & ~new_n2176;
  assign new_n2910 = ~new_n2908 & ~new_n2909;
  assign new_n2911 = ~new_n1794 & ~new_n2910;
  assign new_n2912 = new_n1727 & new_n2911;
  assign new_n2913 = ~new_n2907 & ~new_n2912;
  assign new_n2914 = lo18 & ~new_n1700;
  assign new_n2915 = ~lo18 & new_n2402;
  assign new_n2916 = lo18 & ~new_n2402;
  assign new_n2917 = ~new_n2915 & ~new_n2916;
  assign new_n2918 = lo43 & ~new_n2917;
  assign new_n2919 = new_n1700 & new_n2918;
  assign li18 = new_n2914 | new_n2919;
  assign new_n2921 = new_n2913 & li18;
  assign new_n2922 = ~new_n2913 & ~li18;
  assign new_n2923 = ~new_n2921 & ~new_n2922;
  assign new_n2924 = new_n2906 & new_n2923;
  assign new_n2925 = new_n2889 & new_n2924;
  assign new_n2926 = new_n2850 & new_n2925;
  assign new_n2927 = new_n2767 & new_n2926;
  assign new_n2928 = ~lo12 & ~lo14;
  assign new_n2929 = ~lo10 & new_n2928;
  assign new_n2930 = ~lo11 & new_n2929;
  assign new_n2931 = ~lo13 & new_n2930;
  assign new_n2932 = new_n1722 & ~new_n2931;
  assign new_n2933 = ~new_n2927 & new_n2932;
  assign li12 = new_n1700 & new_n2933;
  assign new_n2935 = li05 & new_n1877;
  assign new_n2936 = ~li05 & ~new_n1877;
  assign new_n2937 = ~new_n2935 & ~new_n2936;
  assign new_n2938 = li04 & new_n1863;
  assign new_n2939 = ~li04 & ~new_n1863;
  assign new_n2940 = ~new_n2938 & ~new_n2939;
  assign new_n2941 = new_n2937 & new_n2940;
  assign new_n2942 = li03 & new_n1849;
  assign new_n2943 = ~li03 & ~new_n1849;
  assign new_n2944 = ~new_n2942 & ~new_n2943;
  assign new_n2945 = li02 & new_n1836;
  assign new_n2946 = ~li02 & ~new_n1836;
  assign new_n2947 = ~new_n2945 & ~new_n2946;
  assign new_n2948 = new_n2944 & new_n2947;
  assign new_n2949 = new_n2941 & new_n2948;
  assign new_n2950 = new_n1828 & ~new_n2949;
  assign li13 = new_n1700 & new_n2950;
  assign new_n2952 = ~new_n1727 & ~new_n1794;
  assign new_n2953 = ~new_n1794 & new_n1797;
  assign new_n2954 = ~new_n1881 & ~new_n2953;
  assign new_n2955 = new_n1727 & ~new_n2954;
  assign new_n2956 = ~new_n2952 & ~new_n2955;
  assign new_n2957 = lo43 & ~new_n1700;
  assign new_n2958 = lo43 & ~li00;
  assign new_n2959 = ~new_n1888 & ~new_n2958;
  assign new_n2960 = new_n1700 & ~new_n2959;
  assign li43 = new_n2957 | new_n2960;
  assign new_n2962 = new_n2956 & li43;
  assign new_n2963 = ~new_n2956 & ~li43;
  assign new_n2964 = ~new_n2962 & ~new_n2963;
  assign new_n2965 = ~lo14 & ~lo15;
  assign new_n2966 = ~lo10 & new_n2965;
  assign new_n2967 = ~lo11 & new_n2966;
  assign new_n2968 = new_n1722 & ~new_n2967;
  assign new_n2969 = ~new_n2964 & new_n2968;
  assign li14 = new_n1700 & new_n2969;
  assign new_n2971 = li00 & new_n1797;
  assign new_n2972 = ~li00 & ~new_n1797;
  assign new_n2973 = ~new_n2971 & ~new_n2972;
  assign new_n2974 = new_n1723 & ~new_n2973;
  assign li15 = new_n1700 & new_n2974;
  assign new_n2976 = li43 & ~new_n2968;
  assign new_n2977 = ~new_n2956 & new_n2968;
  assign li34 = new_n2976 | new_n2977;
  assign new_n2979 = li35 & ~new_n2168;
  assign new_n2980 = ~new_n2154 & new_n2168;
  assign li44 = new_n2979 | new_n2980;
  assign new_n2982 = li36 & ~new_n2168;
  assign new_n2983 = ~new_n2139 & new_n2168;
  assign li45 = new_n2982 | new_n2983;
  assign new_n2985 = li37 & ~new_n2168;
  assign new_n2986 = ~new_n2123 & new_n2168;
  assign li46 = new_n2985 | new_n2986;
  assign new_n2988 = li38 & ~new_n2168;
  assign new_n2989 = ~new_n2108 & new_n2168;
  assign li47 = new_n2988 | new_n2989;
  assign new_n2991 = li39 & ~new_n2168;
  assign new_n2992 = ~new_n2091 & new_n2168;
  assign li48 = new_n2991 | new_n2992;
  assign new_n2994 = li40 & ~new_n2168;
  assign new_n2995 = ~new_n2076 & new_n2168;
  assign li49 = new_n2994 | new_n2995;
  assign new_n2997 = li41 & ~new_n2168;
  assign new_n2998 = ~new_n2060 & new_n2168;
  assign li50 = new_n2997 | new_n2998;
  assign new_n3000 = li42 & ~new_n2168;
  assign new_n3001 = ~new_n2047 & new_n2168;
  assign li51 = new_n3000 | new_n3001;
  assign new_n3003 = li76 & ~new_n2041;
  assign new_n3004 = ~new_n1996 & new_n2041;
  assign li52 = new_n3003 | new_n3004;
  assign new_n3006 = li77 & ~new_n2041;
  assign new_n3007 = ~new_n1981 & new_n2041;
  assign li53 = new_n3006 | new_n3007;
  assign new_n3009 = li78 & ~new_n2041;
  assign new_n3010 = ~new_n1965 & new_n2041;
  assign li54 = new_n3009 | new_n3010;
  assign new_n3012 = li79 & ~new_n2041;
  assign new_n3013 = ~new_n1950 & new_n2041;
  assign li55 = new_n3012 | new_n3013;
  assign new_n3015 = li80 & ~new_n2041;
  assign new_n3016 = ~new_n1933 & new_n2041;
  assign li56 = new_n3015 | new_n3016;
  assign new_n3018 = li81 & ~new_n2041;
  assign new_n3019 = ~new_n1918 & new_n2041;
  assign li57 = new_n3018 | new_n3019;
  assign new_n3021 = li82 & ~new_n2041;
  assign new_n3022 = ~new_n1902 & new_n2041;
  assign li58 = new_n3021 | new_n3022;
  assign new_n3024 = li83 & ~new_n2041;
  assign new_n3025 = ~new_n1886 & new_n2041;
  assign li59 = new_n3024 | new_n3025;
  assign new_n3027 = li18 & ~new_n2932;
  assign new_n3028 = ~new_n2913 & new_n2932;
  assign li60 = new_n3027 | new_n3028;
  assign new_n3030 = li19 & ~new_n2932;
  assign new_n3031 = ~new_n2896 & new_n2932;
  assign li61 = new_n3030 | new_n3031;
  assign new_n3033 = li20 & ~new_n2932;
  assign new_n3034 = ~new_n2878 & new_n2932;
  assign li62 = new_n3033 | new_n3034;
  assign new_n3036 = li21 & ~new_n2932;
  assign new_n3037 = ~new_n2859 & new_n2932;
  assign li63 = new_n3036 | new_n3037;
  assign new_n3039 = li22 & ~new_n2932;
  assign new_n3040 = ~new_n2838 & new_n2932;
  assign li64 = new_n3039 | new_n3040;
  assign new_n3042 = li23 & ~new_n2932;
  assign new_n3043 = ~new_n2819 & new_n2932;
  assign li65 = new_n3042 | new_n3043;
  assign new_n3045 = li24 & ~new_n2932;
  assign new_n3046 = ~new_n2799 & new_n2932;
  assign li66 = new_n3045 | new_n3046;
  assign new_n3048 = li25 & ~new_n2932;
  assign new_n3049 = ~new_n2778 & new_n2932;
  assign li67 = new_n3048 | new_n3049;
  assign new_n3051 = li26 & ~new_n2932;
  assign new_n3052 = ~new_n2754 & new_n2932;
  assign li68 = new_n3051 | new_n3052;
  assign new_n3054 = li27 & ~new_n2932;
  assign new_n3055 = ~new_n2735 & new_n2932;
  assign li69 = new_n3054 | new_n3055;
  assign new_n3057 = li28 & ~new_n2932;
  assign new_n3058 = ~new_n2715 & new_n2932;
  assign li70 = new_n3057 | new_n3058;
  assign new_n3060 = li29 & ~new_n2932;
  assign new_n3061 = ~new_n2694 & new_n2932;
  assign li71 = new_n3060 | new_n3061;
  assign new_n3063 = li30 & ~new_n2932;
  assign new_n3064 = ~new_n2671 & new_n2932;
  assign li72 = new_n3063 | new_n3064;
  assign new_n3066 = li31 & ~new_n2932;
  assign new_n3067 = ~new_n2652 & new_n2932;
  assign li73 = new_n3066 | new_n3067;
  assign new_n3069 = li32 & ~new_n2932;
  assign new_n3070 = ~new_n2632 & new_n2932;
  assign li74 = new_n3069 | new_n3070;
  assign new_n3072 = li33 & ~new_n2932;
  assign new_n3073 = ~new_n2396 & new_n2932;
  assign li75 = new_n3072 | new_n3073;
  assign new_n3075 = lo15 & ~li16;
  assign po0 = ~li17 & new_n3075;
  assign new_n3077 = lo11 & ~li16;
  assign po1 = ~li17 & new_n3077;
  assign new_n3079 = lo14 & ~li16;
  assign po2 = ~li17 & new_n3079;
  assign new_n3081 = lo13 & ~li16;
  assign po3 = ~li17 & new_n3081;
  always @ (posedge clock) begin
    lo00 <= li00;
    lo01 <= li01;
    lo02 <= li02;
    lo03 <= li03;
    lo04 <= li04;
    lo05 <= li05;
    lo06 <= li06;
    lo07 <= li07;
    lo08 <= li08;
    lo09 <= li09;
    lo10 <= li10;
    lo11 <= li11;
    lo12 <= li12;
    lo13 <= li13;
    lo14 <= li14;
    lo15 <= li15;
    lo16 <= li16;
    lo17 <= li17;
    lo18 <= li18;
    lo19 <= li19;
    lo20 <= li20;
    lo21 <= li21;
    lo22 <= li22;
    lo23 <= li23;
    lo24 <= li24;
    lo25 <= li25;
    lo26 <= li26;
    lo27 <= li27;
    lo28 <= li28;
    lo29 <= li29;
    lo30 <= li30;
    lo31 <= li31;
    lo32 <= li32;
    lo33 <= li33;
    lo34 <= li34;
    lo35 <= li35;
    lo36 <= li36;
    lo37 <= li37;
    lo38 <= li38;
    lo39 <= li39;
    lo40 <= li40;
    lo41 <= li41;
    lo42 <= li42;
    lo43 <= li43;
    lo44 <= li44;
    lo45 <= li45;
    lo46 <= li46;
    lo47 <= li47;
    lo48 <= li48;
    lo49 <= li49;
    lo50 <= li50;
    lo51 <= li51;
    lo52 <= li52;
    lo53 <= li53;
    lo54 <= li54;
    lo55 <= li55;
    lo56 <= li56;
    lo57 <= li57;
    lo58 <= li58;
    lo59 <= li59;
    lo60 <= li60;
    lo61 <= li61;
    lo62 <= li62;
    lo63 <= li63;
    lo64 <= li64;
    lo65 <= li65;
    lo66 <= li66;
    lo67 <= li67;
    lo68 <= li68;
    lo69 <= li69;
    lo70 <= li70;
    lo71 <= li71;
    lo72 <= li72;
    lo73 <= li73;
    lo74 <= li74;
    lo75 <= li75;
    lo76 <= li76;
    lo77 <= li77;
    lo78 <= li78;
    lo79 <= li79;
    lo80 <= li80;
    lo81 <= li81;
    lo82 <= li82;
    lo83 <= li83;
  end
  initial begin
    lo00 <= 1'b0;
    lo01 <= 1'b0;
    lo02 <= 1'b0;
    lo03 <= 1'b0;
    lo04 <= 1'b0;
    lo05 <= 1'b0;
    lo06 <= 1'b0;
    lo07 <= 1'b0;
    lo08 <= 1'b0;
    lo09 <= 1'b0;
    lo10 <= 1'b0;
    lo11 <= 1'b0;
    lo12 <= 1'b0;
    lo13 <= 1'b0;
    lo14 <= 1'b0;
    lo15 <= 1'b0;
    lo16 <= 1'b0;
    lo17 <= 1'b0;
    lo18 <= 1'b0;
    lo19 <= 1'b0;
    lo20 <= 1'b0;
    lo21 <= 1'b0;
    lo22 <= 1'b0;
    lo23 <= 1'b0;
    lo24 <= 1'b0;
    lo25 <= 1'b0;
    lo26 <= 1'b0;
    lo27 <= 1'b0;
    lo28 <= 1'b0;
    lo29 <= 1'b0;
    lo30 <= 1'b0;
    lo31 <= 1'b0;
    lo32 <= 1'b0;
    lo33 <= 1'b0;
    lo34 <= 1'b0;
    lo35 <= 1'b0;
    lo36 <= 1'b0;
    lo37 <= 1'b0;
    lo38 <= 1'b0;
    lo39 <= 1'b0;
    lo40 <= 1'b0;
    lo41 <= 1'b0;
    lo42 <= 1'b0;
    lo43 <= 1'b0;
    lo44 <= 1'b0;
    lo45 <= 1'b0;
    lo46 <= 1'b0;
    lo47 <= 1'b0;
    lo48 <= 1'b0;
    lo49 <= 1'b0;
    lo50 <= 1'b0;
    lo51 <= 1'b0;
    lo52 <= 1'b0;
    lo53 <= 1'b0;
    lo54 <= 1'b0;
    lo55 <= 1'b0;
    lo56 <= 1'b0;
    lo57 <= 1'b0;
    lo58 <= 1'b0;
    lo59 <= 1'b0;
    lo60 <= 1'b0;
    lo61 <= 1'b0;
    lo62 <= 1'b0;
    lo63 <= 1'b0;
    lo64 <= 1'b0;
    lo65 <= 1'b0;
    lo66 <= 1'b0;
    lo67 <= 1'b0;
    lo68 <= 1'b0;
    lo69 <= 1'b0;
    lo70 <= 1'b0;
    lo71 <= 1'b0;
    lo72 <= 1'b0;
    lo73 <= 1'b0;
    lo74 <= 1'b0;
    lo75 <= 1'b0;
    lo76 <= 1'b0;
    lo77 <= 1'b0;
    lo78 <= 1'b0;
    lo79 <= 1'b0;
    lo80 <= 1'b0;
    lo81 <= 1'b0;
    lo82 <= 1'b0;
    lo83 <= 1'b0;
  end
endmodule


