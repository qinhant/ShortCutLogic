// Benchmark "fifo" written by ABC on Mon Apr 22 15:24:05 2024

module fifo ( clock, 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14  );
  input  clock;
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14;
  reg lo00, lo01, lo02, lo03, lo04, lo05, lo06, lo07, lo08, lo09, lo10,
    lo11, lo12, lo13, lo14, lo15, lo16, lo17, lo18, lo19, lo20, lo21, lo22,
    lo23, lo24, lo25, lo26, lo27, lo28, lo29, lo30, lo31, lo32, lo33, lo34,
    lo35, lo36, lo37, lo38, lo39, lo40, lo41, lo42, lo43, lo44, lo45, lo46,
    lo47, lo48, lo49, lo50, lo51, lo52, lo53, lo54, lo55, lo56, lo57, lo58,
    lo59, lo60, lo61, lo62, lo63, lo64, lo65, lo66, lo67, lo68, lo69, lo70,
    lo71, lo72, lo73, lo74, lo75, lo76, lo77, lo78, lo79, lo80, lo81, lo82,
    lo83, lo84, lo85, lo86, lo87;
  wire new_n292, new_n293, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n347, new_n348, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n358,
    new_n359, new_n360, new_n361, new_n362, new_n363, new_n364, new_n365,
    new_n366, new_n367, new_n368, new_n369, new_n370, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n397, new_n398, new_n399, new_n400, new_n401, new_n402,
    new_n403, new_n404, new_n405, new_n406, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n418, new_n419, new_n420, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n497,
    new_n498, new_n499, new_n500, new_n501, new_n502, new_n503, new_n504,
    new_n505, new_n506, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n541, new_n542, new_n543, new_n545,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n788, new_n789, new_n791,
    new_n792, new_n794, new_n795, new_n797, new_n798, new_n800, new_n801,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n813, new_n814, new_n816, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n825, new_n826, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n850, new_n851, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n869, new_n870, new_n872, new_n873,
    new_n875, new_n876, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n889, new_n890, new_n892, new_n893,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n911, new_n912, new_n914,
    new_n915, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n939, new_n940, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    li00, li01, li02, li03, li04, li05, li06, li07, li08, li09, li10, li11,
    li12, li13, li14, li15, li16, li17, li18, li19, li20, li21, li22, li23,
    li24, li25, li26, li27, li28, li29, li30, li31, li32, li33, li34, li35,
    li36, li37, li38, li39, li40, li41, li42, li43, li44, li45, li46, li47,
    li48, li49, li50, li51, li52, li53, li54, li55, li56, li57, li58, li59,
    li60, li61, li62, li63, li64, li65, li66, li67, li68, li69, li70, li71,
    li72, li73, li74, li75, li76, li77, li78, li79, li80, li81, li82, li83,
    li84, li85, li86, li87;
  assign new_n292 = ~lo08 & ~lo09;
  assign new_n293 = ~lo10 & new_n292;
  assign po08 = ~lo11 & new_n293;
  assign po09 = lo11 & new_n293;
  assign new_n296 = pi03 & ~po08;
  assign new_n297 = lo00 & ~new_n296;
  assign new_n298 = lo53 & ~lo85;
  assign new_n299 = lo45 & lo85;
  assign new_n300 = ~new_n298 & ~new_n299;
  assign new_n301 = lo87 & ~new_n300;
  assign new_n302 = lo26 & ~lo85;
  assign new_n303 = lo77 & lo85;
  assign new_n304 = ~new_n302 & ~new_n303;
  assign new_n305 = ~lo87 & ~new_n304;
  assign new_n306 = ~new_n301 & ~new_n305;
  assign new_n307 = lo86 & new_n306;
  assign new_n308 = lo69 & ~lo85;
  assign new_n309 = lo61 & lo85;
  assign new_n310 = ~new_n308 & ~new_n309;
  assign new_n311 = lo87 & ~new_n310;
  assign new_n312 = lo18 & ~lo85;
  assign new_n313 = lo34 & lo85;
  assign new_n314 = ~new_n312 & ~new_n313;
  assign new_n315 = ~lo87 & ~new_n314;
  assign new_n316 = ~new_n311 & ~new_n315;
  assign new_n317 = ~lo86 & new_n316;
  assign new_n318 = new_n296 & ~new_n317;
  assign new_n319 = ~new_n307 & new_n318;
  assign new_n320 = ~new_n297 & ~new_n319;
  assign li00 = ~pi00 & ~new_n320;
  assign new_n322 = lo01 & ~new_n296;
  assign new_n323 = lo54 & ~lo85;
  assign new_n324 = lo46 & lo85;
  assign new_n325 = ~new_n323 & ~new_n324;
  assign new_n326 = lo87 & ~new_n325;
  assign new_n327 = lo27 & ~lo85;
  assign new_n328 = lo78 & lo85;
  assign new_n329 = ~new_n327 & ~new_n328;
  assign new_n330 = ~lo87 & ~new_n329;
  assign new_n331 = ~new_n326 & ~new_n330;
  assign new_n332 = lo86 & new_n331;
  assign new_n333 = lo70 & ~lo85;
  assign new_n334 = lo62 & lo85;
  assign new_n335 = ~new_n333 & ~new_n334;
  assign new_n336 = lo87 & ~new_n335;
  assign new_n337 = lo19 & ~lo85;
  assign new_n338 = lo35 & lo85;
  assign new_n339 = ~new_n337 & ~new_n338;
  assign new_n340 = ~lo87 & ~new_n339;
  assign new_n341 = ~new_n336 & ~new_n340;
  assign new_n342 = ~lo86 & new_n341;
  assign new_n343 = new_n296 & ~new_n342;
  assign new_n344 = ~new_n332 & new_n343;
  assign new_n345 = ~new_n322 & ~new_n344;
  assign li01 = ~pi00 & ~new_n345;
  assign new_n347 = lo02 & ~new_n296;
  assign new_n348 = lo55 & ~lo85;
  assign new_n349 = lo47 & lo85;
  assign new_n350 = ~new_n348 & ~new_n349;
  assign new_n351 = lo87 & ~new_n350;
  assign new_n352 = lo28 & ~lo85;
  assign new_n353 = lo79 & lo85;
  assign new_n354 = ~new_n352 & ~new_n353;
  assign new_n355 = ~lo87 & ~new_n354;
  assign new_n356 = ~new_n351 & ~new_n355;
  assign new_n357 = lo86 & new_n356;
  assign new_n358 = lo71 & ~lo85;
  assign new_n359 = lo63 & lo85;
  assign new_n360 = ~new_n358 & ~new_n359;
  assign new_n361 = lo87 & ~new_n360;
  assign new_n362 = lo20 & ~lo85;
  assign new_n363 = lo36 & lo85;
  assign new_n364 = ~new_n362 & ~new_n363;
  assign new_n365 = ~lo87 & ~new_n364;
  assign new_n366 = ~new_n361 & ~new_n365;
  assign new_n367 = ~lo86 & new_n366;
  assign new_n368 = new_n296 & ~new_n367;
  assign new_n369 = ~new_n357 & new_n368;
  assign new_n370 = ~new_n347 & ~new_n369;
  assign li02 = ~pi00 & ~new_n370;
  assign new_n372 = lo03 & ~new_n296;
  assign new_n373 = lo56 & ~lo85;
  assign new_n374 = lo48 & lo85;
  assign new_n375 = ~new_n373 & ~new_n374;
  assign new_n376 = lo87 & ~new_n375;
  assign new_n377 = lo29 & ~lo85;
  assign new_n378 = lo80 & lo85;
  assign new_n379 = ~new_n377 & ~new_n378;
  assign new_n380 = ~lo87 & ~new_n379;
  assign new_n381 = ~new_n376 & ~new_n380;
  assign new_n382 = lo86 & new_n381;
  assign new_n383 = lo72 & ~lo85;
  assign new_n384 = lo64 & lo85;
  assign new_n385 = ~new_n383 & ~new_n384;
  assign new_n386 = lo87 & ~new_n385;
  assign new_n387 = lo21 & ~lo85;
  assign new_n388 = lo37 & lo85;
  assign new_n389 = ~new_n387 & ~new_n388;
  assign new_n390 = ~lo87 & ~new_n389;
  assign new_n391 = ~new_n386 & ~new_n390;
  assign new_n392 = ~lo86 & new_n391;
  assign new_n393 = new_n296 & ~new_n392;
  assign new_n394 = ~new_n382 & new_n393;
  assign new_n395 = ~new_n372 & ~new_n394;
  assign li03 = ~pi00 & ~new_n395;
  assign new_n397 = lo04 & ~new_n296;
  assign new_n398 = lo57 & ~lo85;
  assign new_n399 = lo49 & lo85;
  assign new_n400 = ~new_n398 & ~new_n399;
  assign new_n401 = lo87 & ~new_n400;
  assign new_n402 = lo30 & ~lo85;
  assign new_n403 = lo81 & lo85;
  assign new_n404 = ~new_n402 & ~new_n403;
  assign new_n405 = ~lo87 & ~new_n404;
  assign new_n406 = ~new_n401 & ~new_n405;
  assign new_n407 = lo86 & new_n406;
  assign new_n408 = lo73 & ~lo85;
  assign new_n409 = lo65 & lo85;
  assign new_n410 = ~new_n408 & ~new_n409;
  assign new_n411 = lo87 & ~new_n410;
  assign new_n412 = lo22 & ~lo85;
  assign new_n413 = lo38 & lo85;
  assign new_n414 = ~new_n412 & ~new_n413;
  assign new_n415 = ~lo87 & ~new_n414;
  assign new_n416 = ~new_n411 & ~new_n415;
  assign new_n417 = ~lo86 & new_n416;
  assign new_n418 = new_n296 & ~new_n417;
  assign new_n419 = ~new_n407 & new_n418;
  assign new_n420 = ~new_n397 & ~new_n419;
  assign li04 = ~pi00 & ~new_n420;
  assign new_n422 = lo05 & ~new_n296;
  assign new_n423 = lo58 & ~lo85;
  assign new_n424 = lo50 & lo85;
  assign new_n425 = ~new_n423 & ~new_n424;
  assign new_n426 = lo87 & ~new_n425;
  assign new_n427 = lo31 & ~lo85;
  assign new_n428 = lo82 & lo85;
  assign new_n429 = ~new_n427 & ~new_n428;
  assign new_n430 = ~lo87 & ~new_n429;
  assign new_n431 = ~new_n426 & ~new_n430;
  assign new_n432 = lo86 & new_n431;
  assign new_n433 = lo74 & ~lo85;
  assign new_n434 = lo66 & lo85;
  assign new_n435 = ~new_n433 & ~new_n434;
  assign new_n436 = lo87 & ~new_n435;
  assign new_n437 = lo23 & ~lo85;
  assign new_n438 = lo39 & lo85;
  assign new_n439 = ~new_n437 & ~new_n438;
  assign new_n440 = ~lo87 & ~new_n439;
  assign new_n441 = ~new_n436 & ~new_n440;
  assign new_n442 = ~lo86 & new_n441;
  assign new_n443 = new_n296 & ~new_n442;
  assign new_n444 = ~new_n432 & new_n443;
  assign new_n445 = ~new_n422 & ~new_n444;
  assign li05 = ~pi00 & ~new_n445;
  assign new_n447 = lo06 & ~new_n296;
  assign new_n448 = lo59 & ~lo85;
  assign new_n449 = lo51 & lo85;
  assign new_n450 = ~new_n448 & ~new_n449;
  assign new_n451 = lo87 & ~new_n450;
  assign new_n452 = lo32 & ~lo85;
  assign new_n453 = lo83 & lo85;
  assign new_n454 = ~new_n452 & ~new_n453;
  assign new_n455 = ~lo87 & ~new_n454;
  assign new_n456 = ~new_n451 & ~new_n455;
  assign new_n457 = lo86 & new_n456;
  assign new_n458 = lo75 & ~lo85;
  assign new_n459 = lo67 & lo85;
  assign new_n460 = ~new_n458 & ~new_n459;
  assign new_n461 = lo87 & ~new_n460;
  assign new_n462 = lo24 & ~lo85;
  assign new_n463 = lo40 & lo85;
  assign new_n464 = ~new_n462 & ~new_n463;
  assign new_n465 = ~lo87 & ~new_n464;
  assign new_n466 = ~new_n461 & ~new_n465;
  assign new_n467 = ~lo86 & new_n466;
  assign new_n468 = new_n296 & ~new_n467;
  assign new_n469 = ~new_n457 & new_n468;
  assign new_n470 = ~new_n447 & ~new_n469;
  assign li06 = ~pi00 & ~new_n470;
  assign new_n472 = lo07 & ~new_n296;
  assign new_n473 = lo60 & ~lo85;
  assign new_n474 = lo52 & lo85;
  assign new_n475 = ~new_n473 & ~new_n474;
  assign new_n476 = lo87 & ~new_n475;
  assign new_n477 = lo33 & ~lo85;
  assign new_n478 = lo84 & lo85;
  assign new_n479 = ~new_n477 & ~new_n478;
  assign new_n480 = ~lo87 & ~new_n479;
  assign new_n481 = ~new_n476 & ~new_n480;
  assign new_n482 = lo86 & new_n481;
  assign new_n483 = lo76 & ~lo85;
  assign new_n484 = lo68 & lo85;
  assign new_n485 = ~new_n483 & ~new_n484;
  assign new_n486 = lo87 & ~new_n485;
  assign new_n487 = lo25 & ~lo85;
  assign new_n488 = lo41 & lo85;
  assign new_n489 = ~new_n487 & ~new_n488;
  assign new_n490 = ~lo87 & ~new_n489;
  assign new_n491 = ~new_n486 & ~new_n490;
  assign new_n492 = ~lo86 & new_n491;
  assign new_n493 = new_n296 & ~new_n492;
  assign new_n494 = ~new_n482 & new_n493;
  assign new_n495 = ~new_n472 & ~new_n494;
  assign li07 = ~pi00 & ~new_n495;
  assign new_n497 = pi02 & ~po09;
  assign new_n498 = ~new_n296 & new_n497;
  assign new_n499 = new_n296 & ~new_n497;
  assign new_n500 = ~new_n498 & ~new_n499;
  assign new_n501 = ~lo08 & new_n500;
  assign new_n502 = new_n296 & new_n497;
  assign new_n503 = ~new_n296 & ~new_n497;
  assign new_n504 = ~new_n502 & ~new_n503;
  assign new_n505 = lo08 & new_n504;
  assign new_n506 = ~pi00 & ~new_n505;
  assign li08 = ~new_n501 & new_n506;
  assign new_n508 = ~lo09 & new_n497;
  assign new_n509 = ~pi02 & lo09;
  assign new_n510 = ~new_n508 & ~new_n509;
  assign new_n511 = lo08 & new_n510;
  assign new_n512 = ~lo08 & ~new_n510;
  assign new_n513 = ~new_n511 & ~new_n512;
  assign new_n514 = new_n504 & ~new_n513;
  assign new_n515 = ~lo09 & new_n500;
  assign new_n516 = ~pi00 & ~new_n515;
  assign li09 = ~new_n514 & new_n516;
  assign new_n518 = ~new_n509 & ~new_n511;
  assign new_n519 = pi02 & lo10;
  assign new_n520 = ~lo10 & ~new_n497;
  assign new_n521 = ~new_n519 & ~new_n520;
  assign new_n522 = ~new_n518 & new_n521;
  assign new_n523 = new_n518 & ~new_n521;
  assign new_n524 = ~new_n522 & ~new_n523;
  assign new_n525 = new_n504 & new_n524;
  assign new_n526 = ~lo10 & new_n500;
  assign new_n527 = ~pi00 & ~new_n526;
  assign li10 = ~new_n525 & new_n527;
  assign new_n529 = new_n511 & new_n519;
  assign new_n530 = new_n292 & new_n520;
  assign new_n531 = ~new_n529 & ~new_n530;
  assign new_n532 = new_n504 & ~new_n531;
  assign new_n533 = ~lo11 & ~new_n532;
  assign new_n534 = lo11 & new_n532;
  assign new_n535 = ~pi00 & ~new_n534;
  assign li11 = ~new_n533 & new_n535;
  assign new_n537 = lo12 & new_n296;
  assign new_n538 = ~lo12 & ~new_n296;
  assign new_n539 = ~pi00 & ~new_n538;
  assign li12 = ~new_n537 & new_n539;
  assign new_n541 = lo13 & new_n537;
  assign new_n542 = ~lo13 & ~new_n537;
  assign new_n543 = ~pi00 & ~new_n542;
  assign li13 = ~new_n541 & new_n543;
  assign new_n545 = lo14 & new_n541;
  assign new_n546 = ~lo14 & ~new_n541;
  assign new_n547 = ~pi00 & ~new_n546;
  assign li14 = ~new_n545 & new_n547;
  assign new_n549 = lo15 & new_n497;
  assign new_n550 = ~lo15 & ~new_n497;
  assign new_n551 = ~pi00 & ~new_n550;
  assign li15 = ~new_n549 & new_n551;
  assign new_n553 = lo16 & new_n549;
  assign new_n554 = ~lo16 & ~new_n549;
  assign new_n555 = ~pi00 & ~new_n554;
  assign li16 = ~new_n553 & new_n555;
  assign new_n557 = ~lo17 & ~new_n553;
  assign new_n558 = lo16 & lo17;
  assign new_n559 = new_n549 & new_n558;
  assign new_n560 = ~pi00 & ~new_n559;
  assign li17 = ~new_n557 & new_n560;
  assign new_n562 = ~lo16 & ~lo17;
  assign new_n563 = ~lo15 & new_n562;
  assign new_n564 = ~pi04 & new_n497;
  assign new_n565 = lo34 & ~lo44;
  assign new_n566 = lo44 & lo61;
  assign new_n567 = lo42 & ~new_n566;
  assign new_n568 = ~new_n565 & new_n567;
  assign new_n569 = lo44 & lo69;
  assign new_n570 = lo18 & ~lo44;
  assign new_n571 = ~new_n569 & ~new_n570;
  assign new_n572 = ~lo42 & new_n571;
  assign new_n573 = ~new_n568 & ~new_n572;
  assign new_n574 = ~lo43 & new_n573;
  assign new_n575 = lo44 & lo53;
  assign new_n576 = lo26 & ~lo44;
  assign new_n577 = ~new_n575 & ~new_n576;
  assign new_n578 = ~lo42 & new_n577;
  assign new_n579 = ~lo44 & lo77;
  assign new_n580 = lo44 & lo45;
  assign new_n581 = lo42 & ~new_n580;
  assign new_n582 = ~new_n579 & new_n581;
  assign new_n583 = lo43 & ~new_n582;
  assign new_n584 = ~new_n578 & new_n583;
  assign new_n585 = ~new_n497 & ~new_n584;
  assign new_n586 = ~new_n574 & new_n585;
  assign new_n587 = ~new_n564 & ~new_n586;
  assign new_n588 = new_n563 & new_n587;
  assign new_n589 = lo18 & ~new_n563;
  assign li18 = new_n588 | new_n589;
  assign new_n591 = ~pi05 & new_n497;
  assign new_n592 = lo35 & ~lo44;
  assign new_n593 = lo44 & lo62;
  assign new_n594 = lo42 & ~new_n593;
  assign new_n595 = ~new_n592 & new_n594;
  assign new_n596 = lo44 & lo70;
  assign new_n597 = lo19 & ~lo44;
  assign new_n598 = ~new_n596 & ~new_n597;
  assign new_n599 = ~lo42 & new_n598;
  assign new_n600 = ~new_n595 & ~new_n599;
  assign new_n601 = ~lo43 & new_n600;
  assign new_n602 = lo44 & lo54;
  assign new_n603 = lo27 & ~lo44;
  assign new_n604 = ~new_n602 & ~new_n603;
  assign new_n605 = ~lo42 & new_n604;
  assign new_n606 = ~lo44 & lo78;
  assign new_n607 = lo44 & lo46;
  assign new_n608 = lo42 & ~new_n607;
  assign new_n609 = ~new_n606 & new_n608;
  assign new_n610 = lo43 & ~new_n609;
  assign new_n611 = ~new_n605 & new_n610;
  assign new_n612 = ~new_n497 & ~new_n611;
  assign new_n613 = ~new_n601 & new_n612;
  assign new_n614 = ~new_n591 & ~new_n613;
  assign new_n615 = new_n563 & new_n614;
  assign new_n616 = lo19 & ~new_n563;
  assign li19 = new_n615 | new_n616;
  assign new_n618 = ~pi06 & new_n497;
  assign new_n619 = lo36 & ~lo44;
  assign new_n620 = lo44 & lo63;
  assign new_n621 = lo42 & ~new_n620;
  assign new_n622 = ~new_n619 & new_n621;
  assign new_n623 = lo44 & lo71;
  assign new_n624 = lo20 & ~lo44;
  assign new_n625 = ~new_n623 & ~new_n624;
  assign new_n626 = ~lo42 & new_n625;
  assign new_n627 = ~new_n622 & ~new_n626;
  assign new_n628 = ~lo43 & new_n627;
  assign new_n629 = lo44 & lo55;
  assign new_n630 = lo28 & ~lo44;
  assign new_n631 = ~new_n629 & ~new_n630;
  assign new_n632 = ~lo42 & new_n631;
  assign new_n633 = ~lo44 & lo79;
  assign new_n634 = lo44 & lo47;
  assign new_n635 = lo42 & ~new_n634;
  assign new_n636 = ~new_n633 & new_n635;
  assign new_n637 = lo43 & ~new_n636;
  assign new_n638 = ~new_n632 & new_n637;
  assign new_n639 = ~new_n497 & ~new_n638;
  assign new_n640 = ~new_n628 & new_n639;
  assign new_n641 = ~new_n618 & ~new_n640;
  assign new_n642 = new_n563 & new_n641;
  assign new_n643 = lo20 & ~new_n563;
  assign li20 = new_n642 | new_n643;
  assign new_n645 = ~pi07 & new_n497;
  assign new_n646 = lo37 & ~lo44;
  assign new_n647 = lo44 & lo64;
  assign new_n648 = lo42 & ~new_n647;
  assign new_n649 = ~new_n646 & new_n648;
  assign new_n650 = lo44 & lo72;
  assign new_n651 = lo21 & ~lo44;
  assign new_n652 = ~new_n650 & ~new_n651;
  assign new_n653 = ~lo42 & new_n652;
  assign new_n654 = ~new_n649 & ~new_n653;
  assign new_n655 = ~lo43 & new_n654;
  assign new_n656 = lo44 & lo56;
  assign new_n657 = lo29 & ~lo44;
  assign new_n658 = ~new_n656 & ~new_n657;
  assign new_n659 = ~lo42 & new_n658;
  assign new_n660 = ~lo44 & lo80;
  assign new_n661 = lo44 & lo48;
  assign new_n662 = lo42 & ~new_n661;
  assign new_n663 = ~new_n660 & new_n662;
  assign new_n664 = lo43 & ~new_n663;
  assign new_n665 = ~new_n659 & new_n664;
  assign new_n666 = ~new_n497 & ~new_n665;
  assign new_n667 = ~new_n655 & new_n666;
  assign new_n668 = ~new_n645 & ~new_n667;
  assign new_n669 = new_n563 & new_n668;
  assign new_n670 = lo21 & ~new_n563;
  assign li21 = new_n669 | new_n670;
  assign new_n672 = ~pi08 & new_n497;
  assign new_n673 = lo38 & ~lo44;
  assign new_n674 = lo44 & lo65;
  assign new_n675 = lo42 & ~new_n674;
  assign new_n676 = ~new_n673 & new_n675;
  assign new_n677 = lo44 & lo73;
  assign new_n678 = lo22 & ~lo44;
  assign new_n679 = ~new_n677 & ~new_n678;
  assign new_n680 = ~lo42 & new_n679;
  assign new_n681 = ~new_n676 & ~new_n680;
  assign new_n682 = ~lo43 & new_n681;
  assign new_n683 = lo44 & lo57;
  assign new_n684 = lo30 & ~lo44;
  assign new_n685 = ~new_n683 & ~new_n684;
  assign new_n686 = ~lo42 & new_n685;
  assign new_n687 = ~lo44 & lo81;
  assign new_n688 = lo44 & lo49;
  assign new_n689 = lo42 & ~new_n688;
  assign new_n690 = ~new_n687 & new_n689;
  assign new_n691 = lo43 & ~new_n690;
  assign new_n692 = ~new_n686 & new_n691;
  assign new_n693 = ~new_n497 & ~new_n692;
  assign new_n694 = ~new_n682 & new_n693;
  assign new_n695 = ~new_n672 & ~new_n694;
  assign new_n696 = new_n563 & new_n695;
  assign new_n697 = lo22 & ~new_n563;
  assign li22 = new_n696 | new_n697;
  assign new_n699 = ~pi09 & new_n497;
  assign new_n700 = lo39 & ~lo44;
  assign new_n701 = lo44 & lo66;
  assign new_n702 = lo42 & ~new_n701;
  assign new_n703 = ~new_n700 & new_n702;
  assign new_n704 = lo44 & lo74;
  assign new_n705 = lo23 & ~lo44;
  assign new_n706 = ~new_n704 & ~new_n705;
  assign new_n707 = ~lo42 & new_n706;
  assign new_n708 = ~new_n703 & ~new_n707;
  assign new_n709 = ~lo43 & new_n708;
  assign new_n710 = lo44 & lo58;
  assign new_n711 = lo31 & ~lo44;
  assign new_n712 = ~new_n710 & ~new_n711;
  assign new_n713 = ~lo42 & new_n712;
  assign new_n714 = ~lo44 & lo82;
  assign new_n715 = lo44 & lo50;
  assign new_n716 = lo42 & ~new_n715;
  assign new_n717 = ~new_n714 & new_n716;
  assign new_n718 = lo43 & ~new_n717;
  assign new_n719 = ~new_n713 & new_n718;
  assign new_n720 = ~new_n497 & ~new_n719;
  assign new_n721 = ~new_n709 & new_n720;
  assign new_n722 = ~new_n699 & ~new_n721;
  assign new_n723 = new_n563 & new_n722;
  assign new_n724 = lo23 & ~new_n563;
  assign li23 = new_n723 | new_n724;
  assign new_n726 = ~pi10 & new_n497;
  assign new_n727 = lo40 & ~lo44;
  assign new_n728 = lo44 & lo67;
  assign new_n729 = lo42 & ~new_n728;
  assign new_n730 = ~new_n727 & new_n729;
  assign new_n731 = lo44 & lo75;
  assign new_n732 = lo24 & ~lo44;
  assign new_n733 = ~new_n731 & ~new_n732;
  assign new_n734 = ~lo42 & new_n733;
  assign new_n735 = ~new_n730 & ~new_n734;
  assign new_n736 = ~lo43 & new_n735;
  assign new_n737 = lo44 & lo59;
  assign new_n738 = lo32 & ~lo44;
  assign new_n739 = ~new_n737 & ~new_n738;
  assign new_n740 = ~lo42 & new_n739;
  assign new_n741 = ~lo44 & lo83;
  assign new_n742 = lo44 & lo51;
  assign new_n743 = lo42 & ~new_n742;
  assign new_n744 = ~new_n741 & new_n743;
  assign new_n745 = lo43 & ~new_n744;
  assign new_n746 = ~new_n740 & new_n745;
  assign new_n747 = ~new_n497 & ~new_n746;
  assign new_n748 = ~new_n736 & new_n747;
  assign new_n749 = ~new_n726 & ~new_n748;
  assign new_n750 = new_n563 & new_n749;
  assign new_n751 = lo24 & ~new_n563;
  assign li24 = new_n750 | new_n751;
  assign new_n753 = ~pi11 & new_n497;
  assign new_n754 = lo41 & ~lo44;
  assign new_n755 = lo44 & lo68;
  assign new_n756 = lo42 & ~new_n755;
  assign new_n757 = ~new_n754 & new_n756;
  assign new_n758 = lo44 & lo76;
  assign new_n759 = lo25 & ~lo44;
  assign new_n760 = ~new_n758 & ~new_n759;
  assign new_n761 = ~lo42 & new_n760;
  assign new_n762 = ~new_n757 & ~new_n761;
  assign new_n763 = ~lo43 & new_n762;
  assign new_n764 = lo44 & lo60;
  assign new_n765 = lo33 & ~lo44;
  assign new_n766 = ~new_n764 & ~new_n765;
  assign new_n767 = ~lo42 & new_n766;
  assign new_n768 = ~lo44 & lo84;
  assign new_n769 = lo44 & lo52;
  assign new_n770 = lo42 & ~new_n769;
  assign new_n771 = ~new_n768 & new_n770;
  assign new_n772 = lo43 & ~new_n771;
  assign new_n773 = ~new_n767 & new_n772;
  assign new_n774 = ~new_n497 & ~new_n773;
  assign new_n775 = ~new_n763 & new_n774;
  assign new_n776 = ~new_n753 & ~new_n775;
  assign new_n777 = new_n563 & new_n776;
  assign new_n778 = lo25 & ~new_n563;
  assign li25 = new_n777 | new_n778;
  assign new_n780 = lo16 & ~lo17;
  assign new_n781 = ~lo15 & new_n780;
  assign new_n782 = new_n587 & new_n781;
  assign new_n783 = lo26 & ~new_n781;
  assign li26 = new_n782 | new_n783;
  assign new_n785 = lo27 & ~new_n781;
  assign new_n786 = new_n614 & new_n781;
  assign li27 = new_n785 | new_n786;
  assign new_n788 = lo28 & ~new_n781;
  assign new_n789 = new_n641 & new_n781;
  assign li28 = new_n788 | new_n789;
  assign new_n791 = new_n668 & new_n781;
  assign new_n792 = lo29 & ~new_n781;
  assign li29 = new_n791 | new_n792;
  assign new_n794 = new_n695 & new_n781;
  assign new_n795 = lo30 & ~new_n781;
  assign li30 = new_n794 | new_n795;
  assign new_n797 = lo31 & ~new_n781;
  assign new_n798 = new_n722 & new_n781;
  assign li31 = new_n797 | new_n798;
  assign new_n800 = lo32 & ~new_n781;
  assign new_n801 = new_n749 & new_n781;
  assign li32 = new_n800 | new_n801;
  assign new_n803 = lo33 & ~new_n781;
  assign new_n804 = new_n776 & new_n781;
  assign li33 = new_n803 | new_n804;
  assign new_n806 = lo15 & new_n562;
  assign new_n807 = new_n587 & new_n806;
  assign new_n808 = lo34 & ~new_n806;
  assign li34 = new_n807 | new_n808;
  assign new_n810 = lo35 & ~new_n806;
  assign new_n811 = new_n614 & new_n806;
  assign li35 = new_n810 | new_n811;
  assign new_n813 = lo36 & ~new_n806;
  assign new_n814 = new_n641 & new_n806;
  assign li36 = new_n813 | new_n814;
  assign new_n816 = new_n668 & new_n806;
  assign new_n817 = lo37 & ~new_n806;
  assign li37 = new_n816 | new_n817;
  assign new_n819 = new_n695 & new_n806;
  assign new_n820 = lo38 & ~new_n806;
  assign li38 = new_n819 | new_n820;
  assign new_n822 = lo39 & ~new_n806;
  assign new_n823 = new_n722 & new_n806;
  assign li39 = new_n822 | new_n823;
  assign new_n825 = lo40 & ~new_n806;
  assign new_n826 = new_n749 & new_n806;
  assign li40 = new_n825 | new_n826;
  assign new_n828 = lo41 & ~new_n806;
  assign new_n829 = new_n776 & new_n806;
  assign li41 = new_n828 | new_n829;
  assign new_n831 = lo15 & new_n558;
  assign new_n832 = new_n587 & new_n831;
  assign new_n833 = lo45 & ~new_n831;
  assign li45 = new_n832 | new_n833;
  assign new_n835 = lo46 & ~new_n831;
  assign new_n836 = new_n614 & new_n831;
  assign li46 = new_n835 | new_n836;
  assign new_n838 = lo47 & ~new_n831;
  assign new_n839 = new_n641 & new_n831;
  assign li47 = new_n838 | new_n839;
  assign new_n841 = new_n668 & new_n831;
  assign new_n842 = lo48 & ~new_n831;
  assign li48 = new_n841 | new_n842;
  assign new_n844 = new_n695 & new_n831;
  assign new_n845 = lo49 & ~new_n831;
  assign li49 = new_n844 | new_n845;
  assign new_n847 = lo50 & ~new_n831;
  assign new_n848 = new_n722 & new_n831;
  assign li50 = new_n847 | new_n848;
  assign new_n850 = new_n749 & new_n831;
  assign new_n851 = lo51 & ~new_n831;
  assign li51 = new_n850 | new_n851;
  assign new_n853 = lo52 & ~new_n831;
  assign new_n854 = new_n776 & new_n831;
  assign li52 = new_n853 | new_n854;
  assign new_n856 = ~lo15 & new_n558;
  assign new_n857 = new_n587 & new_n856;
  assign new_n858 = lo53 & ~new_n856;
  assign li53 = new_n857 | new_n858;
  assign new_n860 = lo54 & ~new_n856;
  assign new_n861 = new_n614 & new_n856;
  assign li54 = new_n860 | new_n861;
  assign new_n863 = lo55 & ~new_n856;
  assign new_n864 = new_n641 & new_n856;
  assign li55 = new_n863 | new_n864;
  assign new_n866 = new_n668 & new_n856;
  assign new_n867 = lo56 & ~new_n856;
  assign li56 = new_n866 | new_n867;
  assign new_n869 = new_n695 & new_n856;
  assign new_n870 = lo57 & ~new_n856;
  assign li57 = new_n869 | new_n870;
  assign new_n872 = lo58 & ~new_n856;
  assign new_n873 = new_n722 & new_n856;
  assign li58 = new_n872 | new_n873;
  assign new_n875 = lo59 & ~new_n856;
  assign new_n876 = new_n749 & new_n856;
  assign li59 = new_n875 | new_n876;
  assign new_n878 = lo60 & ~new_n856;
  assign new_n879 = new_n776 & new_n856;
  assign li60 = new_n878 | new_n879;
  assign new_n881 = ~lo16 & lo17;
  assign new_n882 = lo15 & new_n881;
  assign new_n883 = new_n587 & new_n882;
  assign new_n884 = lo61 & ~new_n882;
  assign li61 = new_n883 | new_n884;
  assign new_n886 = lo62 & ~new_n882;
  assign new_n887 = new_n614 & new_n882;
  assign li62 = new_n886 | new_n887;
  assign new_n889 = lo63 & ~new_n882;
  assign new_n890 = new_n641 & new_n882;
  assign li63 = new_n889 | new_n890;
  assign new_n892 = new_n668 & new_n882;
  assign new_n893 = lo64 & ~new_n882;
  assign li64 = new_n892 | new_n893;
  assign new_n895 = new_n695 & new_n882;
  assign new_n896 = lo65 & ~new_n882;
  assign li65 = new_n895 | new_n896;
  assign new_n898 = lo66 & ~new_n882;
  assign new_n899 = new_n722 & new_n882;
  assign li66 = new_n898 | new_n899;
  assign new_n901 = lo67 & ~new_n882;
  assign new_n902 = new_n749 & new_n882;
  assign li67 = new_n901 | new_n902;
  assign new_n904 = lo68 & ~new_n882;
  assign new_n905 = new_n776 & new_n882;
  assign li68 = new_n904 | new_n905;
  assign new_n907 = ~lo15 & new_n881;
  assign new_n908 = new_n587 & new_n907;
  assign new_n909 = lo69 & ~new_n907;
  assign li69 = new_n908 | new_n909;
  assign new_n911 = lo70 & ~new_n907;
  assign new_n912 = new_n614 & new_n907;
  assign li70 = new_n911 | new_n912;
  assign new_n914 = lo71 & ~new_n907;
  assign new_n915 = new_n641 & new_n907;
  assign li71 = new_n914 | new_n915;
  assign new_n917 = new_n668 & new_n907;
  assign new_n918 = lo72 & ~new_n907;
  assign li72 = new_n917 | new_n918;
  assign new_n920 = new_n695 & new_n907;
  assign new_n921 = lo73 & ~new_n907;
  assign li73 = new_n920 | new_n921;
  assign new_n923 = lo74 & ~new_n907;
  assign new_n924 = new_n722 & new_n907;
  assign li74 = new_n923 | new_n924;
  assign new_n926 = lo75 & ~new_n907;
  assign new_n927 = new_n749 & new_n907;
  assign li75 = new_n926 | new_n927;
  assign new_n929 = lo76 & ~new_n907;
  assign new_n930 = new_n776 & new_n907;
  assign li76 = new_n929 | new_n930;
  assign new_n932 = lo15 & new_n780;
  assign new_n933 = new_n587 & new_n932;
  assign new_n934 = lo77 & ~new_n932;
  assign li77 = new_n933 | new_n934;
  assign new_n936 = lo78 & ~new_n932;
  assign new_n937 = new_n614 & new_n932;
  assign li78 = new_n936 | new_n937;
  assign new_n939 = lo79 & ~new_n932;
  assign new_n940 = new_n641 & new_n932;
  assign li79 = new_n939 | new_n940;
  assign new_n942 = new_n668 & new_n932;
  assign new_n943 = lo80 & ~new_n932;
  assign li80 = new_n942 | new_n943;
  assign new_n945 = new_n695 & new_n932;
  assign new_n946 = lo81 & ~new_n932;
  assign li81 = new_n945 | new_n946;
  assign new_n948 = lo82 & ~new_n932;
  assign new_n949 = new_n722 & new_n932;
  assign li82 = new_n948 | new_n949;
  assign new_n951 = lo83 & ~new_n932;
  assign new_n952 = new_n749 & new_n932;
  assign li83 = new_n951 | new_n952;
  assign new_n954 = lo84 & ~new_n932;
  assign new_n955 = new_n776 & new_n932;
  assign li84 = new_n954 | new_n955;
  assign po14 = ~po08;
  assign po00 = lo00;
  assign po01 = lo01;
  assign po02 = lo02;
  assign po03 = lo03;
  assign po04 = lo04;
  assign po05 = lo05;
  assign po06 = lo06;
  assign po07 = lo07;
  assign po10 = lo08;
  assign po11 = lo09;
  assign po12 = lo10;
  assign po13 = lo11;
  assign li42 = li15;
  assign li43 = li16;
  assign li44 = li17;
  assign li85 = li12;
  assign li86 = li13;
  assign li87 = li14;
  always @ (posedge clock) begin
    lo00 <= li00;
    lo01 <= li01;
    lo02 <= li02;
    lo03 <= li03;
    lo04 <= li04;
    lo05 <= li05;
    lo06 <= li06;
    lo07 <= li07;
    lo08 <= li08;
    lo09 <= li09;
    lo10 <= li10;
    lo11 <= li11;
    lo12 <= li12;
    lo13 <= li13;
    lo14 <= li14;
    lo15 <= li15;
    lo16 <= li16;
    lo17 <= li17;
    lo18 <= li18;
    lo19 <= li19;
    lo20 <= li20;
    lo21 <= li21;
    lo22 <= li22;
    lo23 <= li23;
    lo24 <= li24;
    lo25 <= li25;
    lo26 <= li26;
    lo27 <= li27;
    lo28 <= li28;
    lo29 <= li29;
    lo30 <= li30;
    lo31 <= li31;
    lo32 <= li32;
    lo33 <= li33;
    lo34 <= li34;
    lo35 <= li35;
    lo36 <= li36;
    lo37 <= li37;
    lo38 <= li38;
    lo39 <= li39;
    lo40 <= li40;
    lo41 <= li41;
    lo42 <= li42;
    lo43 <= li43;
    lo44 <= li44;
    lo45 <= li45;
    lo46 <= li46;
    lo47 <= li47;
    lo48 <= li48;
    lo49 <= li49;
    lo50 <= li50;
    lo51 <= li51;
    lo52 <= li52;
    lo53 <= li53;
    lo54 <= li54;
    lo55 <= li55;
    lo56 <= li56;
    lo57 <= li57;
    lo58 <= li58;
    lo59 <= li59;
    lo60 <= li60;
    lo61 <= li61;
    lo62 <= li62;
    lo63 <= li63;
    lo64 <= li64;
    lo65 <= li65;
    lo66 <= li66;
    lo67 <= li67;
    lo68 <= li68;
    lo69 <= li69;
    lo70 <= li70;
    lo71 <= li71;
    lo72 <= li72;
    lo73 <= li73;
    lo74 <= li74;
    lo75 <= li75;
    lo76 <= li76;
    lo77 <= li77;
    lo78 <= li78;
    lo79 <= li79;
    lo80 <= li80;
    lo81 <= li81;
    lo82 <= li82;
    lo83 <= li83;
    lo84 <= li84;
    lo85 <= li85;
    lo86 <= li86;
    lo87 <= li87;
  end
  initial begin
    lo00 <= 1'b0;
    lo01 <= 1'b0;
    lo02 <= 1'b0;
    lo03 <= 1'b0;
    lo04 <= 1'b0;
    lo05 <= 1'b0;
    lo06 <= 1'b0;
    lo07 <= 1'b0;
    lo08 <= 1'b0;
    lo09 <= 1'b0;
    lo10 <= 1'b0;
    lo11 <= 1'b0;
    lo12 <= 1'b0;
    lo13 <= 1'b0;
    lo14 <= 1'b0;
    lo15 <= 1'b0;
    lo16 <= 1'b0;
    lo17 <= 1'b0;
    lo18 <= 1'b0;
    lo19 <= 1'b0;
    lo20 <= 1'b0;
    lo21 <= 1'b0;
    lo22 <= 1'b0;
    lo23 <= 1'b0;
    lo24 <= 1'b0;
    lo25 <= 1'b0;
    lo26 <= 1'b0;
    lo27 <= 1'b0;
    lo28 <= 1'b0;
    lo29 <= 1'b0;
    lo30 <= 1'b0;
    lo31 <= 1'b0;
    lo32 <= 1'b0;
    lo33 <= 1'b0;
    lo34 <= 1'b0;
    lo35 <= 1'b0;
    lo36 <= 1'b0;
    lo37 <= 1'b0;
    lo38 <= 1'b0;
    lo39 <= 1'b0;
    lo40 <= 1'b0;
    lo41 <= 1'b0;
    lo42 <= 1'b0;
    lo43 <= 1'b0;
    lo44 <= 1'b0;
    lo45 <= 1'b0;
    lo46 <= 1'b0;
    lo47 <= 1'b0;
    lo48 <= 1'b0;
    lo49 <= 1'b0;
    lo50 <= 1'b0;
    lo51 <= 1'b0;
    lo52 <= 1'b0;
    lo53 <= 1'b0;
    lo54 <= 1'b0;
    lo55 <= 1'b0;
    lo56 <= 1'b0;
    lo57 <= 1'b0;
    lo58 <= 1'b0;
    lo59 <= 1'b0;
    lo60 <= 1'b0;
    lo61 <= 1'b0;
    lo62 <= 1'b0;
    lo63 <= 1'b0;
    lo64 <= 1'b0;
    lo65 <= 1'b0;
    lo66 <= 1'b0;
    lo67 <= 1'b0;
    lo68 <= 1'b0;
    lo69 <= 1'b0;
    lo70 <= 1'b0;
    lo71 <= 1'b0;
    lo72 <= 1'b0;
    lo73 <= 1'b0;
    lo74 <= 1'b0;
    lo75 <= 1'b0;
    lo76 <= 1'b0;
    lo77 <= 1'b0;
    lo78 <= 1'b0;
    lo79 <= 1'b0;
    lo80 <= 1'b0;
    lo81 <= 1'b0;
    lo82 <= 1'b0;
    lo83 <= 1'b0;
    lo84 <= 1'b0;
    lo85 <= 1'b0;
    lo86 <= 1'b0;
    lo87 <= 1'b0;
  end
endmodule


