// Benchmark "fifo" written by ABC on Thu Apr 25 21:52:19 2024

module fifo ( clock, 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    po0  );
  input  clock;
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11;
  output po0;
  reg lo00, lo01, lo02, lo03, lo04, lo05, lo06, lo07, lo08, lo09, lo10,
    lo11, lo12, lo13, lo14, lo15, lo16, lo17, lo18, lo19, lo20, lo21, lo22,
    lo23, lo24, lo25, lo26, lo27, lo28, lo29, lo30, lo31, lo32, lo33, lo34,
    lo35, lo36, lo37, lo38, lo39, lo40, lo41, lo42, lo43, lo44, lo45, lo46,
    lo47, lo48, lo49, lo50, lo51, lo52, lo53, lo54, lo55, lo56, lo57, lo58,
    lo59, lo60, lo61, lo62, lo63, lo64, lo65, lo66, lo67, lo68, lo69, lo70,
    lo71, lo72, lo73, lo74, lo75, lo76, lo77, lo78, lo79, lo80, lo81;
  wire new_n260, new_n261, new_n262, new_n263, new_n264, new_n265, new_n266,
    new_n267, new_n268, new_n269, new_n270, new_n271, new_n272, new_n273,
    new_n274, new_n275, new_n276, new_n277, new_n278, new_n279, new_n280,
    new_n281, new_n282, new_n283, new_n284, new_n285, new_n286, new_n287,
    new_n289, new_n290, new_n291, new_n292, new_n293, new_n294, new_n295,
    new_n296, new_n297, new_n298, new_n299, new_n300, new_n301, new_n302,
    new_n303, new_n304, new_n305, new_n306, new_n307, new_n308, new_n309,
    new_n310, new_n311, new_n312, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n347, new_n348, new_n349, new_n350, new_n351, new_n352, new_n353,
    new_n354, new_n355, new_n356, new_n357, new_n358, new_n359, new_n360,
    new_n361, new_n362, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n444, new_n445, new_n446, new_n447, new_n448,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n462,
    new_n464, new_n465, new_n466, new_n467, new_n468, new_n469, new_n470,
    new_n471, new_n472, new_n473, new_n474, new_n475, new_n476, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n493,
    new_n494, new_n495, new_n496, new_n497, new_n498, new_n499, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n505, new_n506, new_n507,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n526, new_n527, new_n528, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1175, new_n1176, li00, li01,
    li02, li03, li04, li05, li06, li07, li08, li09, li10, li11, li12, li13,
    li14, li15, li16, li17, li18, li19, li20, li21, li22, li23, li24, li25,
    li26, li27, li28, li29, li30, li31, li32, li33, li34, li35, li36, li37,
    li38, li39, li40, li41, li42, li43, li44, li45, li46, li47, li48, li49,
    li50, li51, li52, li53, li54, li55, li56, li57, li58, li59, li60, li61,
    li62, li63, li64, li65, li66, li67, li68, li69, li70, li71, li72, li73,
    li74, li75, li76, li77, li78, li79, li80, li81;
  assign new_n260 = lo12 & lo34;
  assign new_n261 = ~lo12 & lo58;
  assign new_n262 = ~new_n260 & ~new_n261;
  assign new_n263 = lo13 & ~new_n262;
  assign new_n264 = lo12 & lo66;
  assign new_n265 = ~lo12 & lo74;
  assign new_n266 = ~new_n264 & ~new_n265;
  assign new_n267 = ~lo13 & ~new_n266;
  assign new_n268 = ~new_n263 & ~new_n267;
  assign new_n269 = lo14 & ~new_n268;
  assign new_n270 = lo12 & lo26;
  assign new_n271 = ~lo12 & lo18;
  assign new_n272 = ~new_n270 & ~new_n271;
  assign new_n273 = lo13 & ~new_n272;
  assign new_n274 = lo12 & lo42;
  assign new_n275 = ~lo12 & lo50;
  assign new_n276 = ~new_n274 & ~new_n275;
  assign new_n277 = ~lo13 & ~new_n276;
  assign new_n278 = ~new_n273 & ~new_n277;
  assign new_n279 = ~lo14 & ~new_n278;
  assign new_n280 = ~new_n269 & ~new_n279;
  assign new_n281 = ~lo10 & ~lo11;
  assign new_n282 = ~lo08 & ~lo09;
  assign new_n283 = new_n281 & new_n282;
  assign new_n284 = pi03 & ~new_n283;
  assign new_n285 = ~new_n280 & new_n284;
  assign new_n286 = lo00 & ~new_n284;
  assign new_n287 = ~new_n285 & ~new_n286;
  assign li00 = ~pi00 & ~new_n287;
  assign new_n289 = lo12 & lo35;
  assign new_n290 = ~lo12 & lo59;
  assign new_n291 = ~new_n289 & ~new_n290;
  assign new_n292 = lo13 & ~new_n291;
  assign new_n293 = lo12 & lo67;
  assign new_n294 = ~lo12 & lo75;
  assign new_n295 = ~new_n293 & ~new_n294;
  assign new_n296 = ~lo13 & ~new_n295;
  assign new_n297 = ~new_n292 & ~new_n296;
  assign new_n298 = lo14 & ~new_n297;
  assign new_n299 = lo12 & lo27;
  assign new_n300 = ~lo12 & lo19;
  assign new_n301 = ~new_n299 & ~new_n300;
  assign new_n302 = lo13 & ~new_n301;
  assign new_n303 = lo12 & lo43;
  assign new_n304 = ~lo12 & lo51;
  assign new_n305 = ~new_n303 & ~new_n304;
  assign new_n306 = ~lo13 & ~new_n305;
  assign new_n307 = ~new_n302 & ~new_n306;
  assign new_n308 = ~lo14 & ~new_n307;
  assign new_n309 = ~new_n298 & ~new_n308;
  assign new_n310 = new_n284 & ~new_n309;
  assign new_n311 = lo01 & ~new_n284;
  assign new_n312 = ~new_n310 & ~new_n311;
  assign li01 = ~pi00 & ~new_n312;
  assign new_n314 = lo12 & lo36;
  assign new_n315 = ~lo12 & lo60;
  assign new_n316 = ~new_n314 & ~new_n315;
  assign new_n317 = lo13 & ~new_n316;
  assign new_n318 = lo12 & lo68;
  assign new_n319 = ~lo12 & lo76;
  assign new_n320 = ~new_n318 & ~new_n319;
  assign new_n321 = ~lo13 & ~new_n320;
  assign new_n322 = ~new_n317 & ~new_n321;
  assign new_n323 = lo14 & ~new_n322;
  assign new_n324 = lo12 & lo28;
  assign new_n325 = ~lo12 & lo20;
  assign new_n326 = ~new_n324 & ~new_n325;
  assign new_n327 = lo13 & ~new_n326;
  assign new_n328 = lo12 & lo44;
  assign new_n329 = ~lo12 & lo52;
  assign new_n330 = ~new_n328 & ~new_n329;
  assign new_n331 = ~lo13 & ~new_n330;
  assign new_n332 = ~new_n327 & ~new_n331;
  assign new_n333 = ~lo14 & ~new_n332;
  assign new_n334 = ~new_n323 & ~new_n333;
  assign new_n335 = new_n284 & ~new_n334;
  assign new_n336 = lo02 & ~new_n284;
  assign new_n337 = ~new_n335 & ~new_n336;
  assign li02 = ~pi00 & ~new_n337;
  assign new_n339 = lo12 & lo37;
  assign new_n340 = ~lo12 & lo61;
  assign new_n341 = ~new_n339 & ~new_n340;
  assign new_n342 = lo13 & ~new_n341;
  assign new_n343 = lo12 & lo69;
  assign new_n344 = ~lo12 & lo77;
  assign new_n345 = ~new_n343 & ~new_n344;
  assign new_n346 = ~lo13 & ~new_n345;
  assign new_n347 = ~new_n342 & ~new_n346;
  assign new_n348 = lo14 & ~new_n347;
  assign new_n349 = lo12 & lo29;
  assign new_n350 = ~lo12 & lo21;
  assign new_n351 = ~new_n349 & ~new_n350;
  assign new_n352 = lo13 & ~new_n351;
  assign new_n353 = lo12 & lo45;
  assign new_n354 = ~lo12 & lo53;
  assign new_n355 = ~new_n353 & ~new_n354;
  assign new_n356 = ~lo13 & ~new_n355;
  assign new_n357 = ~new_n352 & ~new_n356;
  assign new_n358 = ~lo14 & ~new_n357;
  assign new_n359 = ~new_n348 & ~new_n358;
  assign new_n360 = new_n284 & ~new_n359;
  assign new_n361 = lo03 & ~new_n284;
  assign new_n362 = ~new_n360 & ~new_n361;
  assign li03 = ~pi00 & ~new_n362;
  assign new_n364 = lo12 & lo38;
  assign new_n365 = ~lo12 & lo62;
  assign new_n366 = ~new_n364 & ~new_n365;
  assign new_n367 = lo13 & ~new_n366;
  assign new_n368 = lo12 & lo70;
  assign new_n369 = ~lo12 & lo78;
  assign new_n370 = ~new_n368 & ~new_n369;
  assign new_n371 = ~lo13 & ~new_n370;
  assign new_n372 = ~new_n367 & ~new_n371;
  assign new_n373 = lo14 & ~new_n372;
  assign new_n374 = lo12 & lo30;
  assign new_n375 = ~lo12 & lo22;
  assign new_n376 = ~new_n374 & ~new_n375;
  assign new_n377 = lo13 & ~new_n376;
  assign new_n378 = lo12 & lo46;
  assign new_n379 = ~lo12 & lo54;
  assign new_n380 = ~new_n378 & ~new_n379;
  assign new_n381 = ~lo13 & ~new_n380;
  assign new_n382 = ~new_n377 & ~new_n381;
  assign new_n383 = ~lo14 & ~new_n382;
  assign new_n384 = ~new_n373 & ~new_n383;
  assign new_n385 = new_n284 & ~new_n384;
  assign new_n386 = lo04 & ~new_n284;
  assign new_n387 = ~new_n385 & ~new_n386;
  assign li04 = ~pi00 & ~new_n387;
  assign new_n389 = lo12 & lo39;
  assign new_n390 = ~lo12 & lo63;
  assign new_n391 = ~new_n389 & ~new_n390;
  assign new_n392 = lo13 & ~new_n391;
  assign new_n393 = lo12 & lo71;
  assign new_n394 = ~lo12 & lo79;
  assign new_n395 = ~new_n393 & ~new_n394;
  assign new_n396 = ~lo13 & ~new_n395;
  assign new_n397 = ~new_n392 & ~new_n396;
  assign new_n398 = lo14 & ~new_n397;
  assign new_n399 = lo12 & lo31;
  assign new_n400 = ~lo12 & lo23;
  assign new_n401 = ~new_n399 & ~new_n400;
  assign new_n402 = lo13 & ~new_n401;
  assign new_n403 = lo12 & lo47;
  assign new_n404 = ~lo12 & lo55;
  assign new_n405 = ~new_n403 & ~new_n404;
  assign new_n406 = ~lo13 & ~new_n405;
  assign new_n407 = ~new_n402 & ~new_n406;
  assign new_n408 = ~lo14 & ~new_n407;
  assign new_n409 = ~new_n398 & ~new_n408;
  assign new_n410 = new_n284 & ~new_n409;
  assign new_n411 = lo05 & ~new_n284;
  assign new_n412 = ~new_n410 & ~new_n411;
  assign li05 = ~pi00 & ~new_n412;
  assign new_n414 = lo12 & lo40;
  assign new_n415 = ~lo12 & lo64;
  assign new_n416 = ~new_n414 & ~new_n415;
  assign new_n417 = lo13 & ~new_n416;
  assign new_n418 = lo12 & lo72;
  assign new_n419 = ~lo12 & lo80;
  assign new_n420 = ~new_n418 & ~new_n419;
  assign new_n421 = ~lo13 & ~new_n420;
  assign new_n422 = ~new_n417 & ~new_n421;
  assign new_n423 = lo14 & ~new_n422;
  assign new_n424 = lo12 & lo32;
  assign new_n425 = ~lo12 & lo24;
  assign new_n426 = ~new_n424 & ~new_n425;
  assign new_n427 = lo13 & ~new_n426;
  assign new_n428 = lo12 & lo48;
  assign new_n429 = ~lo12 & lo56;
  assign new_n430 = ~new_n428 & ~new_n429;
  assign new_n431 = ~lo13 & ~new_n430;
  assign new_n432 = ~new_n427 & ~new_n431;
  assign new_n433 = ~lo14 & ~new_n432;
  assign new_n434 = ~new_n423 & ~new_n433;
  assign new_n435 = new_n284 & ~new_n434;
  assign new_n436 = lo06 & ~new_n284;
  assign new_n437 = ~new_n435 & ~new_n436;
  assign li06 = ~pi00 & ~new_n437;
  assign new_n439 = lo12 & lo41;
  assign new_n440 = ~lo12 & lo65;
  assign new_n441 = ~new_n439 & ~new_n440;
  assign new_n442 = lo13 & ~new_n441;
  assign new_n443 = lo12 & lo73;
  assign new_n444 = ~lo12 & lo81;
  assign new_n445 = ~new_n443 & ~new_n444;
  assign new_n446 = ~lo13 & ~new_n445;
  assign new_n447 = ~new_n442 & ~new_n446;
  assign new_n448 = lo14 & ~new_n447;
  assign new_n449 = lo12 & lo33;
  assign new_n450 = ~lo12 & lo25;
  assign new_n451 = ~new_n449 & ~new_n450;
  assign new_n452 = lo13 & ~new_n451;
  assign new_n453 = lo12 & lo49;
  assign new_n454 = ~lo12 & lo57;
  assign new_n455 = ~new_n453 & ~new_n454;
  assign new_n456 = ~lo13 & ~new_n455;
  assign new_n457 = ~new_n452 & ~new_n456;
  assign new_n458 = ~lo14 & ~new_n457;
  assign new_n459 = ~new_n448 & ~new_n458;
  assign new_n460 = new_n284 & ~new_n459;
  assign new_n461 = lo07 & ~new_n284;
  assign new_n462 = ~new_n460 & ~new_n461;
  assign li07 = ~pi00 & ~new_n462;
  assign new_n464 = ~lo10 & lo11;
  assign new_n465 = new_n282 & new_n464;
  assign new_n466 = pi02 & ~new_n465;
  assign new_n467 = new_n284 & new_n466;
  assign new_n468 = lo08 & new_n467;
  assign new_n469 = ~lo08 & new_n466;
  assign new_n470 = ~lo08 & new_n284;
  assign new_n471 = lo08 & ~new_n284;
  assign new_n472 = ~new_n470 & ~new_n471;
  assign new_n473 = ~new_n466 & ~new_n472;
  assign new_n474 = ~new_n469 & ~new_n473;
  assign new_n475 = ~new_n467 & ~new_n474;
  assign new_n476 = ~new_n468 & ~new_n475;
  assign li08 = ~pi00 & ~new_n476;
  assign new_n478 = lo09 & new_n467;
  assign new_n479 = ~lo08 & lo09;
  assign new_n480 = lo08 & ~lo09;
  assign new_n481 = ~new_n479 & ~new_n480;
  assign new_n482 = new_n466 & ~new_n481;
  assign new_n483 = lo08 & lo09;
  assign new_n484 = ~new_n282 & ~new_n483;
  assign new_n485 = new_n284 & ~new_n484;
  assign new_n486 = lo09 & ~new_n284;
  assign new_n487 = ~new_n485 & ~new_n486;
  assign new_n488 = ~new_n466 & ~new_n487;
  assign new_n489 = ~new_n482 & ~new_n488;
  assign new_n490 = ~new_n467 & ~new_n489;
  assign new_n491 = ~new_n478 & ~new_n490;
  assign li09 = ~pi00 & ~new_n491;
  assign new_n493 = lo10 & new_n467;
  assign new_n494 = lo10 & ~new_n483;
  assign new_n495 = ~lo10 & new_n483;
  assign new_n496 = ~new_n494 & ~new_n495;
  assign new_n497 = new_n466 & ~new_n496;
  assign new_n498 = ~lo10 & new_n282;
  assign new_n499 = lo10 & ~new_n282;
  assign new_n500 = ~new_n498 & ~new_n499;
  assign new_n501 = new_n284 & ~new_n500;
  assign new_n502 = lo10 & ~new_n284;
  assign new_n503 = ~new_n501 & ~new_n502;
  assign new_n504 = ~new_n466 & ~new_n503;
  assign new_n505 = ~new_n497 & ~new_n504;
  assign new_n506 = ~new_n467 & ~new_n505;
  assign new_n507 = ~new_n493 & ~new_n506;
  assign li10 = ~pi00 & ~new_n507;
  assign new_n509 = lo11 & new_n467;
  assign new_n510 = lo10 & new_n483;
  assign new_n511 = lo11 & ~new_n510;
  assign new_n512 = ~lo11 & new_n510;
  assign new_n513 = ~new_n511 & ~new_n512;
  assign new_n514 = new_n466 & ~new_n513;
  assign new_n515 = ~lo11 & new_n498;
  assign new_n516 = lo11 & ~new_n498;
  assign new_n517 = ~new_n515 & ~new_n516;
  assign new_n518 = new_n284 & ~new_n517;
  assign new_n519 = lo11 & ~new_n284;
  assign new_n520 = ~new_n518 & ~new_n519;
  assign new_n521 = ~new_n466 & ~new_n520;
  assign new_n522 = ~new_n514 & ~new_n521;
  assign new_n523 = ~new_n467 & ~new_n522;
  assign new_n524 = ~new_n509 & ~new_n523;
  assign li11 = ~pi00 & ~new_n524;
  assign new_n526 = ~lo12 & new_n284;
  assign new_n527 = lo12 & ~new_n284;
  assign new_n528 = ~new_n526 & ~new_n527;
  assign li12 = ~pi00 & ~new_n528;
  assign new_n530 = ~lo12 & lo13;
  assign new_n531 = lo12 & ~lo13;
  assign new_n532 = ~new_n530 & ~new_n531;
  assign new_n533 = new_n284 & ~new_n532;
  assign new_n534 = lo13 & ~new_n284;
  assign new_n535 = ~new_n533 & ~new_n534;
  assign li13 = ~pi00 & ~new_n535;
  assign new_n537 = lo12 & lo13;
  assign new_n538 = lo14 & ~new_n537;
  assign new_n539 = ~lo14 & new_n537;
  assign new_n540 = ~new_n538 & ~new_n539;
  assign new_n541 = new_n284 & ~new_n540;
  assign new_n542 = lo14 & ~new_n284;
  assign new_n543 = ~new_n541 & ~new_n542;
  assign li14 = ~pi00 & ~new_n543;
  assign new_n545 = ~lo15 & new_n466;
  assign new_n546 = lo15 & ~new_n466;
  assign new_n547 = ~new_n545 & ~new_n546;
  assign li15 = ~pi00 & ~new_n547;
  assign new_n549 = ~lo15 & lo16;
  assign new_n550 = lo15 & ~lo16;
  assign new_n551 = ~new_n549 & ~new_n550;
  assign new_n552 = new_n466 & ~new_n551;
  assign new_n553 = lo16 & ~new_n466;
  assign new_n554 = ~new_n552 & ~new_n553;
  assign li16 = ~pi00 & ~new_n554;
  assign new_n556 = lo15 & lo16;
  assign new_n557 = lo17 & ~new_n556;
  assign new_n558 = ~lo17 & new_n556;
  assign new_n559 = ~new_n557 & ~new_n558;
  assign new_n560 = new_n466 & ~new_n559;
  assign new_n561 = lo17 & ~new_n466;
  assign new_n562 = ~new_n560 & ~new_n561;
  assign li17 = ~pi00 & ~new_n562;
  assign new_n564 = new_n553 & ~new_n561;
  assign new_n565 = ~new_n546 & new_n564;
  assign new_n566 = ~new_n466 & new_n565;
  assign new_n567 = lo15 & lo34;
  assign new_n568 = ~lo15 & lo58;
  assign new_n569 = ~new_n567 & ~new_n568;
  assign new_n570 = lo16 & ~new_n569;
  assign new_n571 = lo15 & lo66;
  assign new_n572 = ~lo15 & lo74;
  assign new_n573 = ~new_n571 & ~new_n572;
  assign new_n574 = ~lo16 & ~new_n573;
  assign new_n575 = ~new_n570 & ~new_n574;
  assign new_n576 = lo17 & ~new_n575;
  assign new_n577 = lo15 & lo26;
  assign new_n578 = ~lo15 & lo18;
  assign new_n579 = ~new_n577 & ~new_n578;
  assign new_n580 = lo16 & ~new_n579;
  assign new_n581 = lo15 & lo42;
  assign new_n582 = ~lo15 & lo50;
  assign new_n583 = ~new_n581 & ~new_n582;
  assign new_n584 = ~lo16 & ~new_n583;
  assign new_n585 = ~new_n580 & ~new_n584;
  assign new_n586 = ~lo17 & ~new_n585;
  assign new_n587 = ~new_n576 & ~new_n586;
  assign new_n588 = ~new_n466 & ~new_n587;
  assign new_n589 = new_n566 & new_n588;
  assign new_n590 = lo17 & new_n466;
  assign new_n591 = lo16 & new_n466;
  assign new_n592 = ~new_n590 & new_n591;
  assign new_n593 = lo15 & new_n466;
  assign new_n594 = new_n592 & ~new_n593;
  assign new_n595 = new_n466 & new_n594;
  assign new_n596 = pi04 & new_n466;
  assign new_n597 = new_n595 & new_n596;
  assign new_n598 = lo18 & ~new_n595;
  assign new_n599 = ~new_n597 & ~new_n598;
  assign new_n600 = ~new_n566 & ~new_n599;
  assign li18 = new_n589 | new_n600;
  assign new_n602 = lo15 & lo35;
  assign new_n603 = ~lo15 & lo59;
  assign new_n604 = ~new_n602 & ~new_n603;
  assign new_n605 = lo16 & ~new_n604;
  assign new_n606 = lo15 & lo67;
  assign new_n607 = ~lo15 & lo75;
  assign new_n608 = ~new_n606 & ~new_n607;
  assign new_n609 = ~lo16 & ~new_n608;
  assign new_n610 = ~new_n605 & ~new_n609;
  assign new_n611 = lo17 & ~new_n610;
  assign new_n612 = lo15 & lo27;
  assign new_n613 = ~lo15 & lo19;
  assign new_n614 = ~new_n612 & ~new_n613;
  assign new_n615 = lo16 & ~new_n614;
  assign new_n616 = lo15 & lo43;
  assign new_n617 = ~lo15 & lo51;
  assign new_n618 = ~new_n616 & ~new_n617;
  assign new_n619 = ~lo16 & ~new_n618;
  assign new_n620 = ~new_n615 & ~new_n619;
  assign new_n621 = ~lo17 & ~new_n620;
  assign new_n622 = ~new_n611 & ~new_n621;
  assign new_n623 = ~new_n466 & ~new_n622;
  assign new_n624 = new_n566 & new_n623;
  assign new_n625 = pi05 & new_n466;
  assign new_n626 = new_n595 & new_n625;
  assign new_n627 = lo19 & ~new_n595;
  assign new_n628 = ~new_n626 & ~new_n627;
  assign new_n629 = ~new_n566 & ~new_n628;
  assign li19 = new_n624 | new_n629;
  assign new_n631 = lo15 & lo36;
  assign new_n632 = ~lo15 & lo60;
  assign new_n633 = ~new_n631 & ~new_n632;
  assign new_n634 = lo16 & ~new_n633;
  assign new_n635 = lo15 & lo68;
  assign new_n636 = ~lo15 & lo76;
  assign new_n637 = ~new_n635 & ~new_n636;
  assign new_n638 = ~lo16 & ~new_n637;
  assign new_n639 = ~new_n634 & ~new_n638;
  assign new_n640 = lo17 & ~new_n639;
  assign new_n641 = lo15 & lo28;
  assign new_n642 = ~lo15 & lo20;
  assign new_n643 = ~new_n641 & ~new_n642;
  assign new_n644 = lo16 & ~new_n643;
  assign new_n645 = lo15 & lo44;
  assign new_n646 = ~lo15 & lo52;
  assign new_n647 = ~new_n645 & ~new_n646;
  assign new_n648 = ~lo16 & ~new_n647;
  assign new_n649 = ~new_n644 & ~new_n648;
  assign new_n650 = ~lo17 & ~new_n649;
  assign new_n651 = ~new_n640 & ~new_n650;
  assign new_n652 = ~new_n466 & ~new_n651;
  assign new_n653 = new_n566 & new_n652;
  assign new_n654 = pi06 & new_n466;
  assign new_n655 = new_n595 & new_n654;
  assign new_n656 = lo20 & ~new_n595;
  assign new_n657 = ~new_n655 & ~new_n656;
  assign new_n658 = ~new_n566 & ~new_n657;
  assign li20 = new_n653 | new_n658;
  assign new_n660 = lo15 & lo37;
  assign new_n661 = ~lo15 & lo61;
  assign new_n662 = ~new_n660 & ~new_n661;
  assign new_n663 = lo16 & ~new_n662;
  assign new_n664 = lo15 & lo69;
  assign new_n665 = ~lo15 & lo77;
  assign new_n666 = ~new_n664 & ~new_n665;
  assign new_n667 = ~lo16 & ~new_n666;
  assign new_n668 = ~new_n663 & ~new_n667;
  assign new_n669 = lo17 & ~new_n668;
  assign new_n670 = lo15 & lo29;
  assign new_n671 = ~lo15 & lo21;
  assign new_n672 = ~new_n670 & ~new_n671;
  assign new_n673 = lo16 & ~new_n672;
  assign new_n674 = lo15 & lo45;
  assign new_n675 = ~lo15 & lo53;
  assign new_n676 = ~new_n674 & ~new_n675;
  assign new_n677 = ~lo16 & ~new_n676;
  assign new_n678 = ~new_n673 & ~new_n677;
  assign new_n679 = ~lo17 & ~new_n678;
  assign new_n680 = ~new_n669 & ~new_n679;
  assign new_n681 = ~new_n466 & ~new_n680;
  assign new_n682 = new_n566 & new_n681;
  assign new_n683 = pi07 & new_n466;
  assign new_n684 = new_n595 & new_n683;
  assign new_n685 = lo21 & ~new_n595;
  assign new_n686 = ~new_n684 & ~new_n685;
  assign new_n687 = ~new_n566 & ~new_n686;
  assign li21 = new_n682 | new_n687;
  assign new_n689 = lo15 & lo38;
  assign new_n690 = ~lo15 & lo62;
  assign new_n691 = ~new_n689 & ~new_n690;
  assign new_n692 = lo16 & ~new_n691;
  assign new_n693 = lo15 & lo70;
  assign new_n694 = ~lo15 & lo78;
  assign new_n695 = ~new_n693 & ~new_n694;
  assign new_n696 = ~lo16 & ~new_n695;
  assign new_n697 = ~new_n692 & ~new_n696;
  assign new_n698 = lo17 & ~new_n697;
  assign new_n699 = lo15 & lo30;
  assign new_n700 = ~lo15 & lo22;
  assign new_n701 = ~new_n699 & ~new_n700;
  assign new_n702 = lo16 & ~new_n701;
  assign new_n703 = lo15 & lo46;
  assign new_n704 = ~lo15 & lo54;
  assign new_n705 = ~new_n703 & ~new_n704;
  assign new_n706 = ~lo16 & ~new_n705;
  assign new_n707 = ~new_n702 & ~new_n706;
  assign new_n708 = ~lo17 & ~new_n707;
  assign new_n709 = ~new_n698 & ~new_n708;
  assign new_n710 = ~new_n466 & ~new_n709;
  assign new_n711 = new_n566 & new_n710;
  assign new_n712 = pi08 & new_n466;
  assign new_n713 = new_n595 & new_n712;
  assign new_n714 = lo22 & ~new_n595;
  assign new_n715 = ~new_n713 & ~new_n714;
  assign new_n716 = ~new_n566 & ~new_n715;
  assign li22 = new_n711 | new_n716;
  assign new_n718 = lo15 & lo39;
  assign new_n719 = ~lo15 & lo63;
  assign new_n720 = ~new_n718 & ~new_n719;
  assign new_n721 = lo16 & ~new_n720;
  assign new_n722 = lo15 & lo71;
  assign new_n723 = ~lo15 & lo79;
  assign new_n724 = ~new_n722 & ~new_n723;
  assign new_n725 = ~lo16 & ~new_n724;
  assign new_n726 = ~new_n721 & ~new_n725;
  assign new_n727 = lo17 & ~new_n726;
  assign new_n728 = lo15 & lo31;
  assign new_n729 = ~lo15 & lo23;
  assign new_n730 = ~new_n728 & ~new_n729;
  assign new_n731 = lo16 & ~new_n730;
  assign new_n732 = lo15 & lo47;
  assign new_n733 = ~lo15 & lo55;
  assign new_n734 = ~new_n732 & ~new_n733;
  assign new_n735 = ~lo16 & ~new_n734;
  assign new_n736 = ~new_n731 & ~new_n735;
  assign new_n737 = ~lo17 & ~new_n736;
  assign new_n738 = ~new_n727 & ~new_n737;
  assign new_n739 = ~new_n466 & ~new_n738;
  assign new_n740 = new_n566 & new_n739;
  assign new_n741 = pi09 & new_n466;
  assign new_n742 = new_n595 & new_n741;
  assign new_n743 = lo23 & ~new_n595;
  assign new_n744 = ~new_n742 & ~new_n743;
  assign new_n745 = ~new_n566 & ~new_n744;
  assign li23 = new_n740 | new_n745;
  assign new_n747 = lo15 & lo40;
  assign new_n748 = ~lo15 & lo64;
  assign new_n749 = ~new_n747 & ~new_n748;
  assign new_n750 = lo16 & ~new_n749;
  assign new_n751 = lo15 & lo72;
  assign new_n752 = ~lo15 & lo80;
  assign new_n753 = ~new_n751 & ~new_n752;
  assign new_n754 = ~lo16 & ~new_n753;
  assign new_n755 = ~new_n750 & ~new_n754;
  assign new_n756 = lo17 & ~new_n755;
  assign new_n757 = lo15 & lo32;
  assign new_n758 = ~lo15 & lo24;
  assign new_n759 = ~new_n757 & ~new_n758;
  assign new_n760 = lo16 & ~new_n759;
  assign new_n761 = lo15 & lo48;
  assign new_n762 = ~lo15 & lo56;
  assign new_n763 = ~new_n761 & ~new_n762;
  assign new_n764 = ~lo16 & ~new_n763;
  assign new_n765 = ~new_n760 & ~new_n764;
  assign new_n766 = ~lo17 & ~new_n765;
  assign new_n767 = ~new_n756 & ~new_n766;
  assign new_n768 = ~new_n466 & ~new_n767;
  assign new_n769 = new_n566 & new_n768;
  assign new_n770 = pi10 & new_n466;
  assign new_n771 = new_n595 & new_n770;
  assign new_n772 = lo24 & ~new_n595;
  assign new_n773 = ~new_n771 & ~new_n772;
  assign new_n774 = ~new_n566 & ~new_n773;
  assign li24 = new_n769 | new_n774;
  assign new_n776 = lo15 & lo41;
  assign new_n777 = ~lo15 & lo65;
  assign new_n778 = ~new_n776 & ~new_n777;
  assign new_n779 = lo16 & ~new_n778;
  assign new_n780 = lo15 & lo73;
  assign new_n781 = ~lo15 & lo81;
  assign new_n782 = ~new_n780 & ~new_n781;
  assign new_n783 = ~lo16 & ~new_n782;
  assign new_n784 = ~new_n779 & ~new_n783;
  assign new_n785 = lo17 & ~new_n784;
  assign new_n786 = lo15 & lo33;
  assign new_n787 = ~lo15 & lo25;
  assign new_n788 = ~new_n786 & ~new_n787;
  assign new_n789 = lo16 & ~new_n788;
  assign new_n790 = lo15 & lo49;
  assign new_n791 = ~lo15 & lo57;
  assign new_n792 = ~new_n790 & ~new_n791;
  assign new_n793 = ~lo16 & ~new_n792;
  assign new_n794 = ~new_n789 & ~new_n793;
  assign new_n795 = ~lo17 & ~new_n794;
  assign new_n796 = ~new_n785 & ~new_n795;
  assign new_n797 = ~new_n466 & ~new_n796;
  assign new_n798 = new_n566 & new_n797;
  assign new_n799 = pi11 & new_n466;
  assign new_n800 = new_n595 & new_n799;
  assign new_n801 = lo25 & ~new_n595;
  assign new_n802 = ~new_n800 & ~new_n801;
  assign new_n803 = ~new_n566 & ~new_n802;
  assign li25 = new_n798 | new_n803;
  assign new_n805 = new_n546 & new_n564;
  assign new_n806 = ~new_n466 & new_n805;
  assign new_n807 = new_n588 & new_n806;
  assign new_n808 = new_n592 & new_n593;
  assign new_n809 = new_n466 & new_n808;
  assign new_n810 = new_n596 & new_n809;
  assign new_n811 = lo26 & ~new_n809;
  assign new_n812 = ~new_n810 & ~new_n811;
  assign new_n813 = ~new_n806 & ~new_n812;
  assign li26 = new_n807 | new_n813;
  assign new_n815 = new_n623 & new_n806;
  assign new_n816 = new_n625 & new_n809;
  assign new_n817 = lo27 & ~new_n809;
  assign new_n818 = ~new_n816 & ~new_n817;
  assign new_n819 = ~new_n806 & ~new_n818;
  assign li27 = new_n815 | new_n819;
  assign new_n821 = new_n652 & new_n806;
  assign new_n822 = new_n654 & new_n809;
  assign new_n823 = lo28 & ~new_n809;
  assign new_n824 = ~new_n822 & ~new_n823;
  assign new_n825 = ~new_n806 & ~new_n824;
  assign li28 = new_n821 | new_n825;
  assign new_n827 = new_n681 & new_n806;
  assign new_n828 = new_n683 & new_n809;
  assign new_n829 = lo29 & ~new_n809;
  assign new_n830 = ~new_n828 & ~new_n829;
  assign new_n831 = ~new_n806 & ~new_n830;
  assign li29 = new_n827 | new_n831;
  assign new_n833 = new_n710 & new_n806;
  assign new_n834 = new_n712 & new_n809;
  assign new_n835 = lo30 & ~new_n809;
  assign new_n836 = ~new_n834 & ~new_n835;
  assign new_n837 = ~new_n806 & ~new_n836;
  assign li30 = new_n833 | new_n837;
  assign new_n839 = new_n739 & new_n806;
  assign new_n840 = new_n741 & new_n809;
  assign new_n841 = lo31 & ~new_n809;
  assign new_n842 = ~new_n840 & ~new_n841;
  assign new_n843 = ~new_n806 & ~new_n842;
  assign li31 = new_n839 | new_n843;
  assign new_n845 = new_n768 & new_n806;
  assign new_n846 = new_n770 & new_n809;
  assign new_n847 = lo32 & ~new_n809;
  assign new_n848 = ~new_n846 & ~new_n847;
  assign new_n849 = ~new_n806 & ~new_n848;
  assign li32 = new_n845 | new_n849;
  assign new_n851 = new_n797 & new_n806;
  assign new_n852 = new_n799 & new_n809;
  assign new_n853 = lo33 & ~new_n809;
  assign new_n854 = ~new_n852 & ~new_n853;
  assign new_n855 = ~new_n806 & ~new_n854;
  assign li33 = new_n851 | new_n855;
  assign new_n857 = new_n553 & new_n561;
  assign new_n858 = new_n546 & new_n857;
  assign new_n859 = ~new_n466 & new_n858;
  assign new_n860 = new_n588 & new_n859;
  assign new_n861 = new_n590 & new_n591;
  assign new_n862 = new_n593 & new_n861;
  assign new_n863 = new_n466 & new_n862;
  assign new_n864 = new_n596 & new_n863;
  assign new_n865 = lo34 & ~new_n863;
  assign new_n866 = ~new_n864 & ~new_n865;
  assign new_n867 = ~new_n859 & ~new_n866;
  assign li34 = new_n860 | new_n867;
  assign new_n869 = new_n623 & new_n859;
  assign new_n870 = new_n625 & new_n863;
  assign new_n871 = lo35 & ~new_n863;
  assign new_n872 = ~new_n870 & ~new_n871;
  assign new_n873 = ~new_n859 & ~new_n872;
  assign li35 = new_n869 | new_n873;
  assign new_n875 = new_n652 & new_n859;
  assign new_n876 = new_n654 & new_n863;
  assign new_n877 = lo36 & ~new_n863;
  assign new_n878 = ~new_n876 & ~new_n877;
  assign new_n879 = ~new_n859 & ~new_n878;
  assign li36 = new_n875 | new_n879;
  assign new_n881 = new_n681 & new_n859;
  assign new_n882 = new_n683 & new_n863;
  assign new_n883 = lo37 & ~new_n863;
  assign new_n884 = ~new_n882 & ~new_n883;
  assign new_n885 = ~new_n859 & ~new_n884;
  assign li37 = new_n881 | new_n885;
  assign new_n887 = new_n710 & new_n859;
  assign new_n888 = new_n712 & new_n863;
  assign new_n889 = lo38 & ~new_n863;
  assign new_n890 = ~new_n888 & ~new_n889;
  assign new_n891 = ~new_n859 & ~new_n890;
  assign li38 = new_n887 | new_n891;
  assign new_n893 = new_n739 & new_n859;
  assign new_n894 = new_n741 & new_n863;
  assign new_n895 = lo39 & ~new_n863;
  assign new_n896 = ~new_n894 & ~new_n895;
  assign new_n897 = ~new_n859 & ~new_n896;
  assign li39 = new_n893 | new_n897;
  assign new_n899 = new_n768 & new_n859;
  assign new_n900 = new_n770 & new_n863;
  assign new_n901 = lo40 & ~new_n863;
  assign new_n902 = ~new_n900 & ~new_n901;
  assign new_n903 = ~new_n859 & ~new_n902;
  assign li40 = new_n899 | new_n903;
  assign new_n905 = new_n797 & new_n859;
  assign new_n906 = new_n799 & new_n863;
  assign new_n907 = lo41 & ~new_n863;
  assign new_n908 = ~new_n906 & ~new_n907;
  assign new_n909 = ~new_n859 & ~new_n908;
  assign li41 = new_n905 | new_n909;
  assign new_n911 = ~new_n553 & ~new_n561;
  assign new_n912 = new_n546 & new_n911;
  assign new_n913 = ~new_n466 & new_n912;
  assign new_n914 = new_n588 & new_n913;
  assign new_n915 = ~new_n590 & ~new_n591;
  assign new_n916 = new_n593 & new_n915;
  assign new_n917 = new_n466 & new_n916;
  assign new_n918 = new_n596 & new_n917;
  assign new_n919 = lo42 & ~new_n917;
  assign new_n920 = ~new_n918 & ~new_n919;
  assign new_n921 = ~new_n913 & ~new_n920;
  assign li42 = new_n914 | new_n921;
  assign new_n923 = new_n623 & new_n913;
  assign new_n924 = new_n625 & new_n917;
  assign new_n925 = lo43 & ~new_n917;
  assign new_n926 = ~new_n924 & ~new_n925;
  assign new_n927 = ~new_n913 & ~new_n926;
  assign li43 = new_n923 | new_n927;
  assign new_n929 = new_n652 & new_n913;
  assign new_n930 = new_n654 & new_n917;
  assign new_n931 = lo44 & ~new_n917;
  assign new_n932 = ~new_n930 & ~new_n931;
  assign new_n933 = ~new_n913 & ~new_n932;
  assign li44 = new_n929 | new_n933;
  assign new_n935 = new_n681 & new_n913;
  assign new_n936 = new_n683 & new_n917;
  assign new_n937 = lo45 & ~new_n917;
  assign new_n938 = ~new_n936 & ~new_n937;
  assign new_n939 = ~new_n913 & ~new_n938;
  assign li45 = new_n935 | new_n939;
  assign new_n941 = new_n710 & new_n913;
  assign new_n942 = new_n712 & new_n917;
  assign new_n943 = lo46 & ~new_n917;
  assign new_n944 = ~new_n942 & ~new_n943;
  assign new_n945 = ~new_n913 & ~new_n944;
  assign li46 = new_n941 | new_n945;
  assign new_n947 = new_n739 & new_n913;
  assign new_n948 = new_n741 & new_n917;
  assign new_n949 = lo47 & ~new_n917;
  assign new_n950 = ~new_n948 & ~new_n949;
  assign new_n951 = ~new_n913 & ~new_n950;
  assign li47 = new_n947 | new_n951;
  assign new_n953 = new_n768 & new_n913;
  assign new_n954 = new_n770 & new_n917;
  assign new_n955 = lo48 & ~new_n917;
  assign new_n956 = ~new_n954 & ~new_n955;
  assign new_n957 = ~new_n913 & ~new_n956;
  assign li48 = new_n953 | new_n957;
  assign new_n959 = new_n797 & new_n913;
  assign new_n960 = new_n799 & new_n917;
  assign new_n961 = lo49 & ~new_n917;
  assign new_n962 = ~new_n960 & ~new_n961;
  assign new_n963 = ~new_n913 & ~new_n962;
  assign li49 = new_n959 | new_n963;
  assign new_n965 = ~new_n546 & new_n911;
  assign new_n966 = ~new_n466 & new_n965;
  assign new_n967 = new_n588 & new_n966;
  assign new_n968 = ~new_n593 & new_n915;
  assign new_n969 = new_n466 & new_n968;
  assign new_n970 = new_n596 & new_n969;
  assign new_n971 = lo50 & ~new_n969;
  assign new_n972 = ~new_n970 & ~new_n971;
  assign new_n973 = ~new_n966 & ~new_n972;
  assign li50 = new_n967 | new_n973;
  assign new_n975 = new_n623 & new_n966;
  assign new_n976 = new_n625 & new_n969;
  assign new_n977 = lo51 & ~new_n969;
  assign new_n978 = ~new_n976 & ~new_n977;
  assign new_n979 = ~new_n966 & ~new_n978;
  assign li51 = new_n975 | new_n979;
  assign new_n981 = new_n652 & new_n966;
  assign new_n982 = new_n654 & new_n969;
  assign new_n983 = lo52 & ~new_n969;
  assign new_n984 = ~new_n982 & ~new_n983;
  assign new_n985 = ~new_n966 & ~new_n984;
  assign li52 = new_n981 | new_n985;
  assign new_n987 = new_n681 & new_n966;
  assign new_n988 = new_n683 & new_n969;
  assign new_n989 = lo53 & ~new_n969;
  assign new_n990 = ~new_n988 & ~new_n989;
  assign new_n991 = ~new_n966 & ~new_n990;
  assign li53 = new_n987 | new_n991;
  assign new_n993 = new_n710 & new_n966;
  assign new_n994 = new_n712 & new_n969;
  assign new_n995 = lo54 & ~new_n969;
  assign new_n996 = ~new_n994 & ~new_n995;
  assign new_n997 = ~new_n966 & ~new_n996;
  assign li54 = new_n993 | new_n997;
  assign new_n999 = new_n739 & new_n966;
  assign new_n1000 = new_n741 & new_n969;
  assign new_n1001 = lo55 & ~new_n969;
  assign new_n1002 = ~new_n1000 & ~new_n1001;
  assign new_n1003 = ~new_n966 & ~new_n1002;
  assign li55 = new_n999 | new_n1003;
  assign new_n1005 = new_n768 & new_n966;
  assign new_n1006 = new_n770 & new_n969;
  assign new_n1007 = lo56 & ~new_n969;
  assign new_n1008 = ~new_n1006 & ~new_n1007;
  assign new_n1009 = ~new_n966 & ~new_n1008;
  assign li56 = new_n1005 | new_n1009;
  assign new_n1011 = new_n797 & new_n966;
  assign new_n1012 = new_n799 & new_n969;
  assign new_n1013 = lo57 & ~new_n969;
  assign new_n1014 = ~new_n1012 & ~new_n1013;
  assign new_n1015 = ~new_n966 & ~new_n1014;
  assign li57 = new_n1011 | new_n1015;
  assign new_n1017 = ~new_n546 & new_n857;
  assign new_n1018 = ~new_n466 & new_n1017;
  assign new_n1019 = new_n588 & new_n1018;
  assign new_n1020 = ~new_n593 & new_n861;
  assign new_n1021 = new_n466 & new_n1020;
  assign new_n1022 = new_n596 & new_n1021;
  assign new_n1023 = lo58 & ~new_n1021;
  assign new_n1024 = ~new_n1022 & ~new_n1023;
  assign new_n1025 = ~new_n1018 & ~new_n1024;
  assign li58 = new_n1019 | new_n1025;
  assign new_n1027 = new_n623 & new_n1018;
  assign new_n1028 = new_n625 & new_n1021;
  assign new_n1029 = lo59 & ~new_n1021;
  assign new_n1030 = ~new_n1028 & ~new_n1029;
  assign new_n1031 = ~new_n1018 & ~new_n1030;
  assign li59 = new_n1027 | new_n1031;
  assign new_n1033 = new_n652 & new_n1018;
  assign new_n1034 = new_n654 & new_n1021;
  assign new_n1035 = lo60 & ~new_n1021;
  assign new_n1036 = ~new_n1034 & ~new_n1035;
  assign new_n1037 = ~new_n1018 & ~new_n1036;
  assign li60 = new_n1033 | new_n1037;
  assign new_n1039 = new_n681 & new_n1018;
  assign new_n1040 = new_n683 & new_n1021;
  assign new_n1041 = lo61 & ~new_n1021;
  assign new_n1042 = ~new_n1040 & ~new_n1041;
  assign new_n1043 = ~new_n1018 & ~new_n1042;
  assign li61 = new_n1039 | new_n1043;
  assign new_n1045 = new_n710 & new_n1018;
  assign new_n1046 = new_n712 & new_n1021;
  assign new_n1047 = lo62 & ~new_n1021;
  assign new_n1048 = ~new_n1046 & ~new_n1047;
  assign new_n1049 = ~new_n1018 & ~new_n1048;
  assign li62 = new_n1045 | new_n1049;
  assign new_n1051 = new_n739 & new_n1018;
  assign new_n1052 = new_n741 & new_n1021;
  assign new_n1053 = lo63 & ~new_n1021;
  assign new_n1054 = ~new_n1052 & ~new_n1053;
  assign new_n1055 = ~new_n1018 & ~new_n1054;
  assign li63 = new_n1051 | new_n1055;
  assign new_n1057 = new_n768 & new_n1018;
  assign new_n1058 = new_n770 & new_n1021;
  assign new_n1059 = lo64 & ~new_n1021;
  assign new_n1060 = ~new_n1058 & ~new_n1059;
  assign new_n1061 = ~new_n1018 & ~new_n1060;
  assign li64 = new_n1057 | new_n1061;
  assign new_n1063 = new_n797 & new_n1018;
  assign new_n1064 = new_n799 & new_n1021;
  assign new_n1065 = lo65 & ~new_n1021;
  assign new_n1066 = ~new_n1064 & ~new_n1065;
  assign new_n1067 = ~new_n1018 & ~new_n1066;
  assign li65 = new_n1063 | new_n1067;
  assign new_n1069 = ~new_n553 & new_n561;
  assign new_n1070 = new_n546 & new_n1069;
  assign new_n1071 = ~new_n466 & new_n1070;
  assign new_n1072 = new_n588 & new_n1071;
  assign new_n1073 = new_n590 & ~new_n591;
  assign new_n1074 = new_n593 & new_n1073;
  assign new_n1075 = new_n466 & new_n1074;
  assign new_n1076 = new_n596 & new_n1075;
  assign new_n1077 = lo66 & ~new_n1075;
  assign new_n1078 = ~new_n1076 & ~new_n1077;
  assign new_n1079 = ~new_n1071 & ~new_n1078;
  assign li66 = new_n1072 | new_n1079;
  assign new_n1081 = new_n623 & new_n1071;
  assign new_n1082 = new_n625 & new_n1075;
  assign new_n1083 = lo67 & ~new_n1075;
  assign new_n1084 = ~new_n1082 & ~new_n1083;
  assign new_n1085 = ~new_n1071 & ~new_n1084;
  assign li67 = new_n1081 | new_n1085;
  assign new_n1087 = new_n652 & new_n1071;
  assign new_n1088 = new_n654 & new_n1075;
  assign new_n1089 = lo68 & ~new_n1075;
  assign new_n1090 = ~new_n1088 & ~new_n1089;
  assign new_n1091 = ~new_n1071 & ~new_n1090;
  assign li68 = new_n1087 | new_n1091;
  assign new_n1093 = new_n681 & new_n1071;
  assign new_n1094 = new_n683 & new_n1075;
  assign new_n1095 = lo69 & ~new_n1075;
  assign new_n1096 = ~new_n1094 & ~new_n1095;
  assign new_n1097 = ~new_n1071 & ~new_n1096;
  assign li69 = new_n1093 | new_n1097;
  assign new_n1099 = new_n710 & new_n1071;
  assign new_n1100 = new_n712 & new_n1075;
  assign new_n1101 = lo70 & ~new_n1075;
  assign new_n1102 = ~new_n1100 & ~new_n1101;
  assign new_n1103 = ~new_n1071 & ~new_n1102;
  assign li70 = new_n1099 | new_n1103;
  assign new_n1105 = new_n739 & new_n1071;
  assign new_n1106 = new_n741 & new_n1075;
  assign new_n1107 = lo71 & ~new_n1075;
  assign new_n1108 = ~new_n1106 & ~new_n1107;
  assign new_n1109 = ~new_n1071 & ~new_n1108;
  assign li71 = new_n1105 | new_n1109;
  assign new_n1111 = new_n768 & new_n1071;
  assign new_n1112 = new_n770 & new_n1075;
  assign new_n1113 = lo72 & ~new_n1075;
  assign new_n1114 = ~new_n1112 & ~new_n1113;
  assign new_n1115 = ~new_n1071 & ~new_n1114;
  assign li72 = new_n1111 | new_n1115;
  assign new_n1117 = new_n797 & new_n1071;
  assign new_n1118 = new_n799 & new_n1075;
  assign new_n1119 = lo73 & ~new_n1075;
  assign new_n1120 = ~new_n1118 & ~new_n1119;
  assign new_n1121 = ~new_n1071 & ~new_n1120;
  assign li73 = new_n1117 | new_n1121;
  assign new_n1123 = ~new_n546 & new_n1069;
  assign new_n1124 = ~new_n466 & new_n1123;
  assign new_n1125 = new_n588 & new_n1124;
  assign new_n1126 = ~new_n593 & new_n1073;
  assign new_n1127 = new_n466 & new_n1126;
  assign new_n1128 = new_n596 & new_n1127;
  assign new_n1129 = lo74 & ~new_n1127;
  assign new_n1130 = ~new_n1128 & ~new_n1129;
  assign new_n1131 = ~new_n1124 & ~new_n1130;
  assign li74 = new_n1125 | new_n1131;
  assign new_n1133 = new_n623 & new_n1124;
  assign new_n1134 = new_n625 & new_n1127;
  assign new_n1135 = lo75 & ~new_n1127;
  assign new_n1136 = ~new_n1134 & ~new_n1135;
  assign new_n1137 = ~new_n1124 & ~new_n1136;
  assign li75 = new_n1133 | new_n1137;
  assign new_n1139 = new_n652 & new_n1124;
  assign new_n1140 = new_n654 & new_n1127;
  assign new_n1141 = lo76 & ~new_n1127;
  assign new_n1142 = ~new_n1140 & ~new_n1141;
  assign new_n1143 = ~new_n1124 & ~new_n1142;
  assign li76 = new_n1139 | new_n1143;
  assign new_n1145 = new_n681 & new_n1124;
  assign new_n1146 = new_n683 & new_n1127;
  assign new_n1147 = lo77 & ~new_n1127;
  assign new_n1148 = ~new_n1146 & ~new_n1147;
  assign new_n1149 = ~new_n1124 & ~new_n1148;
  assign li77 = new_n1145 | new_n1149;
  assign new_n1151 = new_n710 & new_n1124;
  assign new_n1152 = new_n712 & new_n1127;
  assign new_n1153 = lo78 & ~new_n1127;
  assign new_n1154 = ~new_n1152 & ~new_n1153;
  assign new_n1155 = ~new_n1124 & ~new_n1154;
  assign li78 = new_n1151 | new_n1155;
  assign new_n1157 = new_n739 & new_n1124;
  assign new_n1158 = new_n741 & new_n1127;
  assign new_n1159 = lo79 & ~new_n1127;
  assign new_n1160 = ~new_n1158 & ~new_n1159;
  assign new_n1161 = ~new_n1124 & ~new_n1160;
  assign li79 = new_n1157 | new_n1161;
  assign new_n1163 = new_n768 & new_n1124;
  assign new_n1164 = new_n770 & new_n1127;
  assign new_n1165 = lo80 & ~new_n1127;
  assign new_n1166 = ~new_n1164 & ~new_n1165;
  assign new_n1167 = ~new_n1124 & ~new_n1166;
  assign li80 = new_n1163 | new_n1167;
  assign new_n1169 = new_n797 & new_n1124;
  assign new_n1170 = new_n799 & new_n1127;
  assign new_n1171 = lo81 & ~new_n1127;
  assign new_n1172 = ~new_n1170 & ~new_n1171;
  assign new_n1173 = ~new_n1124 & ~new_n1172;
  assign li81 = new_n1169 | new_n1173;
  assign new_n1175 = lo10 & lo11;
  assign new_n1176 = ~new_n464 & ~new_n1175;
  assign po0 = ~new_n465 & ~new_n1176;
  always @ (posedge clock) begin
    lo00 <= li00;
    lo01 <= li01;
    lo02 <= li02;
    lo03 <= li03;
    lo04 <= li04;
    lo05 <= li05;
    lo06 <= li06;
    lo07 <= li07;
    lo08 <= li08;
    lo09 <= li09;
    lo10 <= li10;
    lo11 <= li11;
    lo12 <= li12;
    lo13 <= li13;
    lo14 <= li14;
    lo15 <= li15;
    lo16 <= li16;
    lo17 <= li17;
    lo18 <= li18;
    lo19 <= li19;
    lo20 <= li20;
    lo21 <= li21;
    lo22 <= li22;
    lo23 <= li23;
    lo24 <= li24;
    lo25 <= li25;
    lo26 <= li26;
    lo27 <= li27;
    lo28 <= li28;
    lo29 <= li29;
    lo30 <= li30;
    lo31 <= li31;
    lo32 <= li32;
    lo33 <= li33;
    lo34 <= li34;
    lo35 <= li35;
    lo36 <= li36;
    lo37 <= li37;
    lo38 <= li38;
    lo39 <= li39;
    lo40 <= li40;
    lo41 <= li41;
    lo42 <= li42;
    lo43 <= li43;
    lo44 <= li44;
    lo45 <= li45;
    lo46 <= li46;
    lo47 <= li47;
    lo48 <= li48;
    lo49 <= li49;
    lo50 <= li50;
    lo51 <= li51;
    lo52 <= li52;
    lo53 <= li53;
    lo54 <= li54;
    lo55 <= li55;
    lo56 <= li56;
    lo57 <= li57;
    lo58 <= li58;
    lo59 <= li59;
    lo60 <= li60;
    lo61 <= li61;
    lo62 <= li62;
    lo63 <= li63;
    lo64 <= li64;
    lo65 <= li65;
    lo66 <= li66;
    lo67 <= li67;
    lo68 <= li68;
    lo69 <= li69;
    lo70 <= li70;
    lo71 <= li71;
    lo72 <= li72;
    lo73 <= li73;
    lo74 <= li74;
    lo75 <= li75;
    lo76 <= li76;
    lo77 <= li77;
    lo78 <= li78;
    lo79 <= li79;
    lo80 <= li80;
    lo81 <= li81;
  end
  initial begin
    lo00 <= 1'b0;
    lo01 <= 1'b0;
    lo02 <= 1'b0;
    lo03 <= 1'b0;
    lo04 <= 1'b0;
    lo05 <= 1'b0;
    lo06 <= 1'b0;
    lo07 <= 1'b0;
    lo08 <= 1'b0;
    lo09 <= 1'b0;
    lo10 <= 1'b0;
    lo11 <= 1'b0;
    lo12 <= 1'b0;
    lo13 <= 1'b0;
    lo14 <= 1'b0;
    lo15 <= 1'b0;
    lo16 <= 1'b0;
    lo17 <= 1'b0;
    lo18 <= 1'b0;
    lo19 <= 1'b0;
    lo20 <= 1'b0;
    lo21 <= 1'b0;
    lo22 <= 1'b0;
    lo23 <= 1'b0;
    lo24 <= 1'b0;
    lo25 <= 1'b0;
    lo26 <= 1'b0;
    lo27 <= 1'b0;
    lo28 <= 1'b0;
    lo29 <= 1'b0;
    lo30 <= 1'b0;
    lo31 <= 1'b0;
    lo32 <= 1'b0;
    lo33 <= 1'b0;
    lo34 <= 1'b0;
    lo35 <= 1'b0;
    lo36 <= 1'b0;
    lo37 <= 1'b0;
    lo38 <= 1'b0;
    lo39 <= 1'b0;
    lo40 <= 1'b0;
    lo41 <= 1'b0;
    lo42 <= 1'b0;
    lo43 <= 1'b0;
    lo44 <= 1'b0;
    lo45 <= 1'b0;
    lo46 <= 1'b0;
    lo47 <= 1'b0;
    lo48 <= 1'b0;
    lo49 <= 1'b0;
    lo50 <= 1'b0;
    lo51 <= 1'b0;
    lo52 <= 1'b0;
    lo53 <= 1'b0;
    lo54 <= 1'b0;
    lo55 <= 1'b0;
    lo56 <= 1'b0;
    lo57 <= 1'b0;
    lo58 <= 1'b0;
    lo59 <= 1'b0;
    lo60 <= 1'b0;
    lo61 <= 1'b0;
    lo62 <= 1'b0;
    lo63 <= 1'b0;
    lo64 <= 1'b0;
    lo65 <= 1'b0;
    lo66 <= 1'b0;
    lo67 <= 1'b0;
    lo68 <= 1'b0;
    lo69 <= 1'b0;
    lo70 <= 1'b0;
    lo71 <= 1'b0;
    lo72 <= 1'b0;
    lo73 <= 1'b0;
    lo74 <= 1'b0;
    lo75 <= 1'b0;
    lo76 <= 1'b0;
    lo77 <= 1'b0;
    lo78 <= 1'b0;
    lo79 <= 1'b0;
    lo80 <= 1'b0;
    lo81 <= 1'b0;
  end
endmodule


